module bch_ibm(syndrome1, syndrome2, syndrome3, syndrome4, syndrome5, locator0, locator1, locator2, locator3);
  input [9:0] syndrome1;
  input [9:0] syndrome2;
  input [9:0] syndrome3;
  input [9:0] syndrome4;
  input [9:0] syndrome5;
  output [9:0] locator0;
  output [9:0] locator1;
  output [9:0] locator2;
  output [9:0] locator3;

  wire [9:0] nu0_0;
  wire [9:0] nu0_1;
  wire [9:0] nu0_2;
  wire [9:0] nu0_3;
  wire [9:0] nu2_0;
  wire [9:0] nu2_1;
  wire [9:0] nu2_2;
  wire [9:0] nu2_3;
  wire [9:0] nu4_0;
  wire [9:0] nu4_1;
  wire [9:0] nu4_2;
  wire [9:0] nu4_3;
  wire [9:0] nu6_0;
  wire [9:0] nu6_1;
  wire [9:0] nu6_2;
  wire [9:0] nu6_3;
  wire [9:0] kappa0_0;
  wire [9:0] kappa0_1;
  wire [9:0] kappa0_2;
  wire [9:0] kappa0_3;
  wire [9:0] kappa2_0;
  wire [9:0] kappa2_1;
  wire [9:0] kappa2_2;
  wire [9:0] kappa2_3;
  wire [9:0] kappa4_0;
  wire [9:0] kappa4_1;
  wire [9:0] kappa4_2;
  wire [9:0] kappa4_3;
  wire [9:0] kappa6_0;
  wire [9:0] kappa6_1;
  wire [9:0] kappa6_2;
  wire [9:0] kappa6_3;
  wire [9:0] delta0;
  wire [9:0] delta2;
  wire [9:0] delta4;
  wire [9:0] d0;
  wire [9:0] d2;
  wire [9:0] d4;
  wire [9:0] delta0_x_nu2_0;
  wire [9:0] delta0_x_nu2_1;
  wire [9:0] delta0_x_nu2_2;
  wire [9:0] delta0_x_nu2_3;
  wire [9:0] delta2_x_nu4_0;
  wire [9:0] delta2_x_nu4_1;
  wire [9:0] delta2_x_nu4_2;
  wire [9:0] delta2_x_nu4_3;
  wire [9:0] d0_x_kappa0_0;
  wire [9:0] d0_x_kappa0_1;
  wire [9:0] d0_x_kappa0_2;
  wire [9:0] d0_x_kappa0_3;
  wire [9:0] d2_x_kappa2_0;
  wire [9:0] d2_x_kappa2_1;
  wire [9:0] d2_x_kappa2_2;
  wire [9:0] d2_x_kappa2_3;
  wire [9:0] d4_x_kappa4_0;
  wire [9:0] d4_x_kappa4_1;
  wire [9:0] d4_x_kappa4_2;
  wire [9:0] d4_x_kappa4_3;
  wire [9:0] nu0_0_x_syndrome1;
  wire [9:0] nu2_0_x_syndrome3;
  wire [9:0] nu2_1_x_syndrome2;
  wire [9:0] nu2_2_x_syndrome1;
  wire [9:0] nu4_0_x_syndrome5;
  wire [9:0] nu4_1_x_syndrome4;
  wire [9:0] nu4_2_x_syndrome3;
  wire [9:0] nu4_3_x_syndrome2;
  wire cond0;
  wire cond2;
  wire cond4;

  gfmult gfm_delta0_x_nu2_0(delta0, nu2_0, delta0_x_nu2_0);
  gfmult gfm_delta0_x_nu2_1(delta0, nu2_1, delta0_x_nu2_1);
  gfmult gfm_delta0_x_nu2_2(delta0, nu2_2, delta0_x_nu2_2);
  gfmult gfm_delta0_x_nu2_3(delta0, nu2_3, delta0_x_nu2_3);
  gfmult gfm_delta2_x_nu4_0(delta2, nu4_0, delta2_x_nu4_0);
  gfmult gfm_delta2_x_nu4_1(delta2, nu4_1, delta2_x_nu4_1);
  gfmult gfm_delta2_x_nu4_2(delta2, nu4_2, delta2_x_nu4_2);
  gfmult gfm_delta2_x_nu4_3(delta2, nu4_3, delta2_x_nu4_3);
  gfmult gfm_d0_x_kappa0_0(d0, kappa0_0, d0_x_kappa0_0);
  gfmult gfm_d0_x_kappa0_1(d0, kappa0_1, d0_x_kappa0_1);
  gfmult gfm_d0_x_kappa0_2(d0, kappa0_2, d0_x_kappa0_2);
  gfmult gfm_d0_x_kappa0_3(d0, kappa0_3, d0_x_kappa0_3);
  gfmult gfm_d2_x_kappa2_0(d2, kappa2_0, d2_x_kappa2_0);
  gfmult gfm_d2_x_kappa2_1(d2, kappa2_1, d2_x_kappa2_1);
  gfmult gfm_d2_x_kappa2_2(d2, kappa2_2, d2_x_kappa2_2);
  gfmult gfm_d2_x_kappa2_3(d2, kappa2_3, d2_x_kappa2_3);
  gfmult gfm_d4_x_kappa4_0(d4, kappa4_0, d4_x_kappa4_0);
  gfmult gfm_d4_x_kappa4_1(d4, kappa4_1, d4_x_kappa4_1);
  gfmult gfm_d4_x_kappa4_2(d4, kappa4_2, d4_x_kappa4_2);
  gfmult gfm_d4_x_kappa4_3(d4, kappa4_3, d4_x_kappa4_3);
  gfmult gfm_nu0_0_x_syndrome1(nu0_0, syndrome1, nu0_0_x_syndrome1);
  gfmult gfm_nu2_0_x_syndrome3(nu2_0, syndrome3, nu2_0_x_syndrome3);
  gfmult gfm_nu2_1_x_syndrome2(nu2_1, syndrome2, nu2_1_x_syndrome2);
  gfmult gfm_nu2_2_x_syndrome1(nu2_2, syndrome1, nu2_2_x_syndrome1);
  gfmult gfm_nu4_0_x_syndrome5(nu4_0, syndrome5, nu4_0_x_syndrome5);
  gfmult gfm_nu4_1_x_syndrome4(nu4_1, syndrome4, nu4_1_x_syndrome4);
  gfmult gfm_nu4_2_x_syndrome3(nu4_2, syndrome3, nu4_2_x_syndrome3);
  gfmult gfm_nu4_3_x_syndrome2(nu4_3, syndrome2, nu4_3_x_syndrome2);

  assign locator0 = nu6_0;
  assign locator1 = nu6_1;
  assign locator2 = nu6_2;
  assign locator3 = nu6_3;
  assign nu0_0 = 10'b0000000001;
  assign nu0_1 = 10'b0;
  assign nu0_2 = 10'b0;
  assign nu0_3 = 10'b0;
  assign nu2_0 = nu0_0;
  assign nu2_1 = nu0_1 ^ d0_x_kappa0_0;
  assign nu2_2 = nu0_2 ^ d0_x_kappa0_1;
  assign nu2_3 = nu0_3 ^ d0_x_kappa0_2;
  assign nu4_0 = delta0_x_nu2_0;
  assign nu4_1 = delta0_x_nu2_1 ^ d2_x_kappa2_0;
  assign nu4_2 = delta0_x_nu2_2 ^ d2_x_kappa2_1;
  assign nu4_3 = delta0_x_nu2_3 ^ d2_x_kappa2_2;
  assign nu6_0 = delta2_x_nu4_0;
  assign nu6_1 = delta2_x_nu4_1 ^ d4_x_kappa4_0;
  assign nu6_2 = delta2_x_nu4_2 ^ d4_x_kappa4_1;
  assign nu6_3 = delta2_x_nu4_3 ^ d4_x_kappa4_2;
  assign kappa0_0 = 10'b0000000001;
  assign kappa0_1 = 10'b0;
  assign kappa0_2 = 10'b0;
  assign kappa0_3 = 10'b0;
  assign kappa2_0 = cond0 ? 10'b0 : 10'b0;
  assign kappa2_1 = cond0 ? 10'b0 : nu0_0;
  assign kappa2_2 = cond0 ? kappa0_0 : nu0_1;
  assign kappa2_3 = cond0 ? kappa0_1 : nu0_2;
  assign kappa4_0 = cond2 ? 10'b0 : 10'b0;
  assign kappa4_1 = cond2 ? 10'b0 : nu2_0;
  assign kappa4_2 = cond2 ? kappa2_0 : nu2_1;
  assign kappa4_3 = cond2 ? kappa2_1 : nu2_2;
  assign kappa6_0 = cond4 ? 10'b0 : 10'b0;
  assign kappa6_1 = cond4 ? 10'b0 : nu4_0;
  assign kappa6_2 = cond4 ? kappa4_0 : nu4_1;
  assign kappa6_3 = cond4 ? kappa4_1 : nu4_2;
  assign delta0 = cond0 ? 10'b0000000001 : d0;
  assign delta2 = cond2 ? delta0 : d2;
  assign delta4 = cond4 ? delta2 : d4;
  assign d0 = nu0_0_x_syndrome1 ^ nu0_1;
  assign d2 = nu2_0_x_syndrome3 ^ nu2_1_x_syndrome2 ^ nu2_2_x_syndrome1 ^ nu2_3;
  assign d4 = nu4_0_x_syndrome5 ^ nu4_1_x_syndrome4 ^ nu4_2_x_syndrome3 ^ nu4_3_x_syndrome2;
  assign cond0 = (~| d0) | (| nu0_1) | (| nu0_2) | (| nu0_3);
  assign cond2 = (~| d2) | (| nu2_2) | (| nu2_3);
  assign cond4 = (~| d4) | (| nu4_3);
endmodule
