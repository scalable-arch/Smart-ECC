module bch_chien(received, locator0, locator1, locator2, locator3, codeword);
  input [541:0] received;
  input [9:0] locator0;
  input [9:0] locator1;
  input [9:0] locator2;
  input [9:0] locator3;
  output [541:0] codeword;

  wire [541:0] error;
  wire [9:0] alpha0_0_x_locator0;
  wire [9:0] alpha0_1_x_locator1;
  wire [9:0] alpha0_2_x_locator2;
  wire [9:0] alpha0_3_x_locator3;
  wire [9:0] alpha1_0_x_locator0;
  wire [9:0] alpha1_1_x_locator1;
  wire [9:0] alpha1_2_x_locator2;
  wire [9:0] alpha1_3_x_locator3;
  wire [9:0] alpha2_0_x_locator0;
  wire [9:0] alpha2_1_x_locator1;
  wire [9:0] alpha2_2_x_locator2;
  wire [9:0] alpha2_3_x_locator3;
  wire [9:0] alpha3_0_x_locator0;
  wire [9:0] alpha3_1_x_locator1;
  wire [9:0] alpha3_2_x_locator2;
  wire [9:0] alpha3_3_x_locator3;
  wire [9:0] alpha4_0_x_locator0;
  wire [9:0] alpha4_1_x_locator1;
  wire [9:0] alpha4_2_x_locator2;
  wire [9:0] alpha4_3_x_locator3;
  wire [9:0] alpha5_0_x_locator0;
  wire [9:0] alpha5_1_x_locator1;
  wire [9:0] alpha5_2_x_locator2;
  wire [9:0] alpha5_3_x_locator3;
  wire [9:0] alpha6_0_x_locator0;
  wire [9:0] alpha6_1_x_locator1;
  wire [9:0] alpha6_2_x_locator2;
  wire [9:0] alpha6_3_x_locator3;
  wire [9:0] alpha7_0_x_locator0;
  wire [9:0] alpha7_1_x_locator1;
  wire [9:0] alpha7_2_x_locator2;
  wire [9:0] alpha7_3_x_locator3;
  wire [9:0] alpha8_0_x_locator0;
  wire [9:0] alpha8_1_x_locator1;
  wire [9:0] alpha8_2_x_locator2;
  wire [9:0] alpha8_3_x_locator3;
  wire [9:0] alpha9_0_x_locator0;
  wire [9:0] alpha9_1_x_locator1;
  wire [9:0] alpha9_2_x_locator2;
  wire [9:0] alpha9_3_x_locator3;
  wire [9:0] alpha10_0_x_locator0;
  wire [9:0] alpha10_1_x_locator1;
  wire [9:0] alpha10_2_x_locator2;
  wire [9:0] alpha10_3_x_locator3;
  wire [9:0] alpha11_0_x_locator0;
  wire [9:0] alpha11_1_x_locator1;
  wire [9:0] alpha11_2_x_locator2;
  wire [9:0] alpha11_3_x_locator3;
  wire [9:0] alpha12_0_x_locator0;
  wire [9:0] alpha12_1_x_locator1;
  wire [9:0] alpha12_2_x_locator2;
  wire [9:0] alpha12_3_x_locator3;
  wire [9:0] alpha13_0_x_locator0;
  wire [9:0] alpha13_1_x_locator1;
  wire [9:0] alpha13_2_x_locator2;
  wire [9:0] alpha13_3_x_locator3;
  wire [9:0] alpha14_0_x_locator0;
  wire [9:0] alpha14_1_x_locator1;
  wire [9:0] alpha14_2_x_locator2;
  wire [9:0] alpha14_3_x_locator3;
  wire [9:0] alpha15_0_x_locator0;
  wire [9:0] alpha15_1_x_locator1;
  wire [9:0] alpha15_2_x_locator2;
  wire [9:0] alpha15_3_x_locator3;
  wire [9:0] alpha16_0_x_locator0;
  wire [9:0] alpha16_1_x_locator1;
  wire [9:0] alpha16_2_x_locator2;
  wire [9:0] alpha16_3_x_locator3;
  wire [9:0] alpha17_0_x_locator0;
  wire [9:0] alpha17_1_x_locator1;
  wire [9:0] alpha17_2_x_locator2;
  wire [9:0] alpha17_3_x_locator3;
  wire [9:0] alpha18_0_x_locator0;
  wire [9:0] alpha18_1_x_locator1;
  wire [9:0] alpha18_2_x_locator2;
  wire [9:0] alpha18_3_x_locator3;
  wire [9:0] alpha19_0_x_locator0;
  wire [9:0] alpha19_1_x_locator1;
  wire [9:0] alpha19_2_x_locator2;
  wire [9:0] alpha19_3_x_locator3;
  wire [9:0] alpha20_0_x_locator0;
  wire [9:0] alpha20_1_x_locator1;
  wire [9:0] alpha20_2_x_locator2;
  wire [9:0] alpha20_3_x_locator3;
  wire [9:0] alpha21_0_x_locator0;
  wire [9:0] alpha21_1_x_locator1;
  wire [9:0] alpha21_2_x_locator2;
  wire [9:0] alpha21_3_x_locator3;
  wire [9:0] alpha22_0_x_locator0;
  wire [9:0] alpha22_1_x_locator1;
  wire [9:0] alpha22_2_x_locator2;
  wire [9:0] alpha22_3_x_locator3;
  wire [9:0] alpha23_0_x_locator0;
  wire [9:0] alpha23_1_x_locator1;
  wire [9:0] alpha23_2_x_locator2;
  wire [9:0] alpha23_3_x_locator3;
  wire [9:0] alpha24_0_x_locator0;
  wire [9:0] alpha24_1_x_locator1;
  wire [9:0] alpha24_2_x_locator2;
  wire [9:0] alpha24_3_x_locator3;
  wire [9:0] alpha25_0_x_locator0;
  wire [9:0] alpha25_1_x_locator1;
  wire [9:0] alpha25_2_x_locator2;
  wire [9:0] alpha25_3_x_locator3;
  wire [9:0] alpha26_0_x_locator0;
  wire [9:0] alpha26_1_x_locator1;
  wire [9:0] alpha26_2_x_locator2;
  wire [9:0] alpha26_3_x_locator3;
  wire [9:0] alpha27_0_x_locator0;
  wire [9:0] alpha27_1_x_locator1;
  wire [9:0] alpha27_2_x_locator2;
  wire [9:0] alpha27_3_x_locator3;
  wire [9:0] alpha28_0_x_locator0;
  wire [9:0] alpha28_1_x_locator1;
  wire [9:0] alpha28_2_x_locator2;
  wire [9:0] alpha28_3_x_locator3;
  wire [9:0] alpha29_0_x_locator0;
  wire [9:0] alpha29_1_x_locator1;
  wire [9:0] alpha29_2_x_locator2;
  wire [9:0] alpha29_3_x_locator3;
  wire [9:0] alpha30_0_x_locator0;
  wire [9:0] alpha30_1_x_locator1;
  wire [9:0] alpha30_2_x_locator2;
  wire [9:0] alpha30_3_x_locator3;
  wire [9:0] alpha31_0_x_locator0;
  wire [9:0] alpha31_1_x_locator1;
  wire [9:0] alpha31_2_x_locator2;
  wire [9:0] alpha31_3_x_locator3;
  wire [9:0] alpha32_0_x_locator0;
  wire [9:0] alpha32_1_x_locator1;
  wire [9:0] alpha32_2_x_locator2;
  wire [9:0] alpha32_3_x_locator3;
  wire [9:0] alpha33_0_x_locator0;
  wire [9:0] alpha33_1_x_locator1;
  wire [9:0] alpha33_2_x_locator2;
  wire [9:0] alpha33_3_x_locator3;
  wire [9:0] alpha34_0_x_locator0;
  wire [9:0] alpha34_1_x_locator1;
  wire [9:0] alpha34_2_x_locator2;
  wire [9:0] alpha34_3_x_locator3;
  wire [9:0] alpha35_0_x_locator0;
  wire [9:0] alpha35_1_x_locator1;
  wire [9:0] alpha35_2_x_locator2;
  wire [9:0] alpha35_3_x_locator3;
  wire [9:0] alpha36_0_x_locator0;
  wire [9:0] alpha36_1_x_locator1;
  wire [9:0] alpha36_2_x_locator2;
  wire [9:0] alpha36_3_x_locator3;
  wire [9:0] alpha37_0_x_locator0;
  wire [9:0] alpha37_1_x_locator1;
  wire [9:0] alpha37_2_x_locator2;
  wire [9:0] alpha37_3_x_locator3;
  wire [9:0] alpha38_0_x_locator0;
  wire [9:0] alpha38_1_x_locator1;
  wire [9:0] alpha38_2_x_locator2;
  wire [9:0] alpha38_3_x_locator3;
  wire [9:0] alpha39_0_x_locator0;
  wire [9:0] alpha39_1_x_locator1;
  wire [9:0] alpha39_2_x_locator2;
  wire [9:0] alpha39_3_x_locator3;
  wire [9:0] alpha40_0_x_locator0;
  wire [9:0] alpha40_1_x_locator1;
  wire [9:0] alpha40_2_x_locator2;
  wire [9:0] alpha40_3_x_locator3;
  wire [9:0] alpha41_0_x_locator0;
  wire [9:0] alpha41_1_x_locator1;
  wire [9:0] alpha41_2_x_locator2;
  wire [9:0] alpha41_3_x_locator3;
  wire [9:0] alpha42_0_x_locator0;
  wire [9:0] alpha42_1_x_locator1;
  wire [9:0] alpha42_2_x_locator2;
  wire [9:0] alpha42_3_x_locator3;
  wire [9:0] alpha43_0_x_locator0;
  wire [9:0] alpha43_1_x_locator1;
  wire [9:0] alpha43_2_x_locator2;
  wire [9:0] alpha43_3_x_locator3;
  wire [9:0] alpha44_0_x_locator0;
  wire [9:0] alpha44_1_x_locator1;
  wire [9:0] alpha44_2_x_locator2;
  wire [9:0] alpha44_3_x_locator3;
  wire [9:0] alpha45_0_x_locator0;
  wire [9:0] alpha45_1_x_locator1;
  wire [9:0] alpha45_2_x_locator2;
  wire [9:0] alpha45_3_x_locator3;
  wire [9:0] alpha46_0_x_locator0;
  wire [9:0] alpha46_1_x_locator1;
  wire [9:0] alpha46_2_x_locator2;
  wire [9:0] alpha46_3_x_locator3;
  wire [9:0] alpha47_0_x_locator0;
  wire [9:0] alpha47_1_x_locator1;
  wire [9:0] alpha47_2_x_locator2;
  wire [9:0] alpha47_3_x_locator3;
  wire [9:0] alpha48_0_x_locator0;
  wire [9:0] alpha48_1_x_locator1;
  wire [9:0] alpha48_2_x_locator2;
  wire [9:0] alpha48_3_x_locator3;
  wire [9:0] alpha49_0_x_locator0;
  wire [9:0] alpha49_1_x_locator1;
  wire [9:0] alpha49_2_x_locator2;
  wire [9:0] alpha49_3_x_locator3;
  wire [9:0] alpha50_0_x_locator0;
  wire [9:0] alpha50_1_x_locator1;
  wire [9:0] alpha50_2_x_locator2;
  wire [9:0] alpha50_3_x_locator3;
  wire [9:0] alpha51_0_x_locator0;
  wire [9:0] alpha51_1_x_locator1;
  wire [9:0] alpha51_2_x_locator2;
  wire [9:0] alpha51_3_x_locator3;
  wire [9:0] alpha52_0_x_locator0;
  wire [9:0] alpha52_1_x_locator1;
  wire [9:0] alpha52_2_x_locator2;
  wire [9:0] alpha52_3_x_locator3;
  wire [9:0] alpha53_0_x_locator0;
  wire [9:0] alpha53_1_x_locator1;
  wire [9:0] alpha53_2_x_locator2;
  wire [9:0] alpha53_3_x_locator3;
  wire [9:0] alpha54_0_x_locator0;
  wire [9:0] alpha54_1_x_locator1;
  wire [9:0] alpha54_2_x_locator2;
  wire [9:0] alpha54_3_x_locator3;
  wire [9:0] alpha55_0_x_locator0;
  wire [9:0] alpha55_1_x_locator1;
  wire [9:0] alpha55_2_x_locator2;
  wire [9:0] alpha55_3_x_locator3;
  wire [9:0] alpha56_0_x_locator0;
  wire [9:0] alpha56_1_x_locator1;
  wire [9:0] alpha56_2_x_locator2;
  wire [9:0] alpha56_3_x_locator3;
  wire [9:0] alpha57_0_x_locator0;
  wire [9:0] alpha57_1_x_locator1;
  wire [9:0] alpha57_2_x_locator2;
  wire [9:0] alpha57_3_x_locator3;
  wire [9:0] alpha58_0_x_locator0;
  wire [9:0] alpha58_1_x_locator1;
  wire [9:0] alpha58_2_x_locator2;
  wire [9:0] alpha58_3_x_locator3;
  wire [9:0] alpha59_0_x_locator0;
  wire [9:0] alpha59_1_x_locator1;
  wire [9:0] alpha59_2_x_locator2;
  wire [9:0] alpha59_3_x_locator3;
  wire [9:0] alpha60_0_x_locator0;
  wire [9:0] alpha60_1_x_locator1;
  wire [9:0] alpha60_2_x_locator2;
  wire [9:0] alpha60_3_x_locator3;
  wire [9:0] alpha61_0_x_locator0;
  wire [9:0] alpha61_1_x_locator1;
  wire [9:0] alpha61_2_x_locator2;
  wire [9:0] alpha61_3_x_locator3;
  wire [9:0] alpha62_0_x_locator0;
  wire [9:0] alpha62_1_x_locator1;
  wire [9:0] alpha62_2_x_locator2;
  wire [9:0] alpha62_3_x_locator3;
  wire [9:0] alpha63_0_x_locator0;
  wire [9:0] alpha63_1_x_locator1;
  wire [9:0] alpha63_2_x_locator2;
  wire [9:0] alpha63_3_x_locator3;
  wire [9:0] alpha64_0_x_locator0;
  wire [9:0] alpha64_1_x_locator1;
  wire [9:0] alpha64_2_x_locator2;
  wire [9:0] alpha64_3_x_locator3;
  wire [9:0] alpha65_0_x_locator0;
  wire [9:0] alpha65_1_x_locator1;
  wire [9:0] alpha65_2_x_locator2;
  wire [9:0] alpha65_3_x_locator3;
  wire [9:0] alpha66_0_x_locator0;
  wire [9:0] alpha66_1_x_locator1;
  wire [9:0] alpha66_2_x_locator2;
  wire [9:0] alpha66_3_x_locator3;
  wire [9:0] alpha67_0_x_locator0;
  wire [9:0] alpha67_1_x_locator1;
  wire [9:0] alpha67_2_x_locator2;
  wire [9:0] alpha67_3_x_locator3;
  wire [9:0] alpha68_0_x_locator0;
  wire [9:0] alpha68_1_x_locator1;
  wire [9:0] alpha68_2_x_locator2;
  wire [9:0] alpha68_3_x_locator3;
  wire [9:0] alpha69_0_x_locator0;
  wire [9:0] alpha69_1_x_locator1;
  wire [9:0] alpha69_2_x_locator2;
  wire [9:0] alpha69_3_x_locator3;
  wire [9:0] alpha70_0_x_locator0;
  wire [9:0] alpha70_1_x_locator1;
  wire [9:0] alpha70_2_x_locator2;
  wire [9:0] alpha70_3_x_locator3;
  wire [9:0] alpha71_0_x_locator0;
  wire [9:0] alpha71_1_x_locator1;
  wire [9:0] alpha71_2_x_locator2;
  wire [9:0] alpha71_3_x_locator3;
  wire [9:0] alpha72_0_x_locator0;
  wire [9:0] alpha72_1_x_locator1;
  wire [9:0] alpha72_2_x_locator2;
  wire [9:0] alpha72_3_x_locator3;
  wire [9:0] alpha73_0_x_locator0;
  wire [9:0] alpha73_1_x_locator1;
  wire [9:0] alpha73_2_x_locator2;
  wire [9:0] alpha73_3_x_locator3;
  wire [9:0] alpha74_0_x_locator0;
  wire [9:0] alpha74_1_x_locator1;
  wire [9:0] alpha74_2_x_locator2;
  wire [9:0] alpha74_3_x_locator3;
  wire [9:0] alpha75_0_x_locator0;
  wire [9:0] alpha75_1_x_locator1;
  wire [9:0] alpha75_2_x_locator2;
  wire [9:0] alpha75_3_x_locator3;
  wire [9:0] alpha76_0_x_locator0;
  wire [9:0] alpha76_1_x_locator1;
  wire [9:0] alpha76_2_x_locator2;
  wire [9:0] alpha76_3_x_locator3;
  wire [9:0] alpha77_0_x_locator0;
  wire [9:0] alpha77_1_x_locator1;
  wire [9:0] alpha77_2_x_locator2;
  wire [9:0] alpha77_3_x_locator3;
  wire [9:0] alpha78_0_x_locator0;
  wire [9:0] alpha78_1_x_locator1;
  wire [9:0] alpha78_2_x_locator2;
  wire [9:0] alpha78_3_x_locator3;
  wire [9:0] alpha79_0_x_locator0;
  wire [9:0] alpha79_1_x_locator1;
  wire [9:0] alpha79_2_x_locator2;
  wire [9:0] alpha79_3_x_locator3;
  wire [9:0] alpha80_0_x_locator0;
  wire [9:0] alpha80_1_x_locator1;
  wire [9:0] alpha80_2_x_locator2;
  wire [9:0] alpha80_3_x_locator3;
  wire [9:0] alpha81_0_x_locator0;
  wire [9:0] alpha81_1_x_locator1;
  wire [9:0] alpha81_2_x_locator2;
  wire [9:0] alpha81_3_x_locator3;
  wire [9:0] alpha82_0_x_locator0;
  wire [9:0] alpha82_1_x_locator1;
  wire [9:0] alpha82_2_x_locator2;
  wire [9:0] alpha82_3_x_locator3;
  wire [9:0] alpha83_0_x_locator0;
  wire [9:0] alpha83_1_x_locator1;
  wire [9:0] alpha83_2_x_locator2;
  wire [9:0] alpha83_3_x_locator3;
  wire [9:0] alpha84_0_x_locator0;
  wire [9:0] alpha84_1_x_locator1;
  wire [9:0] alpha84_2_x_locator2;
  wire [9:0] alpha84_3_x_locator3;
  wire [9:0] alpha85_0_x_locator0;
  wire [9:0] alpha85_1_x_locator1;
  wire [9:0] alpha85_2_x_locator2;
  wire [9:0] alpha85_3_x_locator3;
  wire [9:0] alpha86_0_x_locator0;
  wire [9:0] alpha86_1_x_locator1;
  wire [9:0] alpha86_2_x_locator2;
  wire [9:0] alpha86_3_x_locator3;
  wire [9:0] alpha87_0_x_locator0;
  wire [9:0] alpha87_1_x_locator1;
  wire [9:0] alpha87_2_x_locator2;
  wire [9:0] alpha87_3_x_locator3;
  wire [9:0] alpha88_0_x_locator0;
  wire [9:0] alpha88_1_x_locator1;
  wire [9:0] alpha88_2_x_locator2;
  wire [9:0] alpha88_3_x_locator3;
  wire [9:0] alpha89_0_x_locator0;
  wire [9:0] alpha89_1_x_locator1;
  wire [9:0] alpha89_2_x_locator2;
  wire [9:0] alpha89_3_x_locator3;
  wire [9:0] alpha90_0_x_locator0;
  wire [9:0] alpha90_1_x_locator1;
  wire [9:0] alpha90_2_x_locator2;
  wire [9:0] alpha90_3_x_locator3;
  wire [9:0] alpha91_0_x_locator0;
  wire [9:0] alpha91_1_x_locator1;
  wire [9:0] alpha91_2_x_locator2;
  wire [9:0] alpha91_3_x_locator3;
  wire [9:0] alpha92_0_x_locator0;
  wire [9:0] alpha92_1_x_locator1;
  wire [9:0] alpha92_2_x_locator2;
  wire [9:0] alpha92_3_x_locator3;
  wire [9:0] alpha93_0_x_locator0;
  wire [9:0] alpha93_1_x_locator1;
  wire [9:0] alpha93_2_x_locator2;
  wire [9:0] alpha93_3_x_locator3;
  wire [9:0] alpha94_0_x_locator0;
  wire [9:0] alpha94_1_x_locator1;
  wire [9:0] alpha94_2_x_locator2;
  wire [9:0] alpha94_3_x_locator3;
  wire [9:0] alpha95_0_x_locator0;
  wire [9:0] alpha95_1_x_locator1;
  wire [9:0] alpha95_2_x_locator2;
  wire [9:0] alpha95_3_x_locator3;
  wire [9:0] alpha96_0_x_locator0;
  wire [9:0] alpha96_1_x_locator1;
  wire [9:0] alpha96_2_x_locator2;
  wire [9:0] alpha96_3_x_locator3;
  wire [9:0] alpha97_0_x_locator0;
  wire [9:0] alpha97_1_x_locator1;
  wire [9:0] alpha97_2_x_locator2;
  wire [9:0] alpha97_3_x_locator3;
  wire [9:0] alpha98_0_x_locator0;
  wire [9:0] alpha98_1_x_locator1;
  wire [9:0] alpha98_2_x_locator2;
  wire [9:0] alpha98_3_x_locator3;
  wire [9:0] alpha99_0_x_locator0;
  wire [9:0] alpha99_1_x_locator1;
  wire [9:0] alpha99_2_x_locator2;
  wire [9:0] alpha99_3_x_locator3;
  wire [9:0] alpha100_0_x_locator0;
  wire [9:0] alpha100_1_x_locator1;
  wire [9:0] alpha100_2_x_locator2;
  wire [9:0] alpha100_3_x_locator3;
  wire [9:0] alpha101_0_x_locator0;
  wire [9:0] alpha101_1_x_locator1;
  wire [9:0] alpha101_2_x_locator2;
  wire [9:0] alpha101_3_x_locator3;
  wire [9:0] alpha102_0_x_locator0;
  wire [9:0] alpha102_1_x_locator1;
  wire [9:0] alpha102_2_x_locator2;
  wire [9:0] alpha102_3_x_locator3;
  wire [9:0] alpha103_0_x_locator0;
  wire [9:0] alpha103_1_x_locator1;
  wire [9:0] alpha103_2_x_locator2;
  wire [9:0] alpha103_3_x_locator3;
  wire [9:0] alpha104_0_x_locator0;
  wire [9:0] alpha104_1_x_locator1;
  wire [9:0] alpha104_2_x_locator2;
  wire [9:0] alpha104_3_x_locator3;
  wire [9:0] alpha105_0_x_locator0;
  wire [9:0] alpha105_1_x_locator1;
  wire [9:0] alpha105_2_x_locator2;
  wire [9:0] alpha105_3_x_locator3;
  wire [9:0] alpha106_0_x_locator0;
  wire [9:0] alpha106_1_x_locator1;
  wire [9:0] alpha106_2_x_locator2;
  wire [9:0] alpha106_3_x_locator3;
  wire [9:0] alpha107_0_x_locator0;
  wire [9:0] alpha107_1_x_locator1;
  wire [9:0] alpha107_2_x_locator2;
  wire [9:0] alpha107_3_x_locator3;
  wire [9:0] alpha108_0_x_locator0;
  wire [9:0] alpha108_1_x_locator1;
  wire [9:0] alpha108_2_x_locator2;
  wire [9:0] alpha108_3_x_locator3;
  wire [9:0] alpha109_0_x_locator0;
  wire [9:0] alpha109_1_x_locator1;
  wire [9:0] alpha109_2_x_locator2;
  wire [9:0] alpha109_3_x_locator3;
  wire [9:0] alpha110_0_x_locator0;
  wire [9:0] alpha110_1_x_locator1;
  wire [9:0] alpha110_2_x_locator2;
  wire [9:0] alpha110_3_x_locator3;
  wire [9:0] alpha111_0_x_locator0;
  wire [9:0] alpha111_1_x_locator1;
  wire [9:0] alpha111_2_x_locator2;
  wire [9:0] alpha111_3_x_locator3;
  wire [9:0] alpha112_0_x_locator0;
  wire [9:0] alpha112_1_x_locator1;
  wire [9:0] alpha112_2_x_locator2;
  wire [9:0] alpha112_3_x_locator3;
  wire [9:0] alpha113_0_x_locator0;
  wire [9:0] alpha113_1_x_locator1;
  wire [9:0] alpha113_2_x_locator2;
  wire [9:0] alpha113_3_x_locator3;
  wire [9:0] alpha114_0_x_locator0;
  wire [9:0] alpha114_1_x_locator1;
  wire [9:0] alpha114_2_x_locator2;
  wire [9:0] alpha114_3_x_locator3;
  wire [9:0] alpha115_0_x_locator0;
  wire [9:0] alpha115_1_x_locator1;
  wire [9:0] alpha115_2_x_locator2;
  wire [9:0] alpha115_3_x_locator3;
  wire [9:0] alpha116_0_x_locator0;
  wire [9:0] alpha116_1_x_locator1;
  wire [9:0] alpha116_2_x_locator2;
  wire [9:0] alpha116_3_x_locator3;
  wire [9:0] alpha117_0_x_locator0;
  wire [9:0] alpha117_1_x_locator1;
  wire [9:0] alpha117_2_x_locator2;
  wire [9:0] alpha117_3_x_locator3;
  wire [9:0] alpha118_0_x_locator0;
  wire [9:0] alpha118_1_x_locator1;
  wire [9:0] alpha118_2_x_locator2;
  wire [9:0] alpha118_3_x_locator3;
  wire [9:0] alpha119_0_x_locator0;
  wire [9:0] alpha119_1_x_locator1;
  wire [9:0] alpha119_2_x_locator2;
  wire [9:0] alpha119_3_x_locator3;
  wire [9:0] alpha120_0_x_locator0;
  wire [9:0] alpha120_1_x_locator1;
  wire [9:0] alpha120_2_x_locator2;
  wire [9:0] alpha120_3_x_locator3;
  wire [9:0] alpha121_0_x_locator0;
  wire [9:0] alpha121_1_x_locator1;
  wire [9:0] alpha121_2_x_locator2;
  wire [9:0] alpha121_3_x_locator3;
  wire [9:0] alpha122_0_x_locator0;
  wire [9:0] alpha122_1_x_locator1;
  wire [9:0] alpha122_2_x_locator2;
  wire [9:0] alpha122_3_x_locator3;
  wire [9:0] alpha123_0_x_locator0;
  wire [9:0] alpha123_1_x_locator1;
  wire [9:0] alpha123_2_x_locator2;
  wire [9:0] alpha123_3_x_locator3;
  wire [9:0] alpha124_0_x_locator0;
  wire [9:0] alpha124_1_x_locator1;
  wire [9:0] alpha124_2_x_locator2;
  wire [9:0] alpha124_3_x_locator3;
  wire [9:0] alpha125_0_x_locator0;
  wire [9:0] alpha125_1_x_locator1;
  wire [9:0] alpha125_2_x_locator2;
  wire [9:0] alpha125_3_x_locator3;
  wire [9:0] alpha126_0_x_locator0;
  wire [9:0] alpha126_1_x_locator1;
  wire [9:0] alpha126_2_x_locator2;
  wire [9:0] alpha126_3_x_locator3;
  wire [9:0] alpha127_0_x_locator0;
  wire [9:0] alpha127_1_x_locator1;
  wire [9:0] alpha127_2_x_locator2;
  wire [9:0] alpha127_3_x_locator3;
  wire [9:0] alpha128_0_x_locator0;
  wire [9:0] alpha128_1_x_locator1;
  wire [9:0] alpha128_2_x_locator2;
  wire [9:0] alpha128_3_x_locator3;
  wire [9:0] alpha129_0_x_locator0;
  wire [9:0] alpha129_1_x_locator1;
  wire [9:0] alpha129_2_x_locator2;
  wire [9:0] alpha129_3_x_locator3;
  wire [9:0] alpha130_0_x_locator0;
  wire [9:0] alpha130_1_x_locator1;
  wire [9:0] alpha130_2_x_locator2;
  wire [9:0] alpha130_3_x_locator3;
  wire [9:0] alpha131_0_x_locator0;
  wire [9:0] alpha131_1_x_locator1;
  wire [9:0] alpha131_2_x_locator2;
  wire [9:0] alpha131_3_x_locator3;
  wire [9:0] alpha132_0_x_locator0;
  wire [9:0] alpha132_1_x_locator1;
  wire [9:0] alpha132_2_x_locator2;
  wire [9:0] alpha132_3_x_locator3;
  wire [9:0] alpha133_0_x_locator0;
  wire [9:0] alpha133_1_x_locator1;
  wire [9:0] alpha133_2_x_locator2;
  wire [9:0] alpha133_3_x_locator3;
  wire [9:0] alpha134_0_x_locator0;
  wire [9:0] alpha134_1_x_locator1;
  wire [9:0] alpha134_2_x_locator2;
  wire [9:0] alpha134_3_x_locator3;
  wire [9:0] alpha135_0_x_locator0;
  wire [9:0] alpha135_1_x_locator1;
  wire [9:0] alpha135_2_x_locator2;
  wire [9:0] alpha135_3_x_locator3;
  wire [9:0] alpha136_0_x_locator0;
  wire [9:0] alpha136_1_x_locator1;
  wire [9:0] alpha136_2_x_locator2;
  wire [9:0] alpha136_3_x_locator3;
  wire [9:0] alpha137_0_x_locator0;
  wire [9:0] alpha137_1_x_locator1;
  wire [9:0] alpha137_2_x_locator2;
  wire [9:0] alpha137_3_x_locator3;
  wire [9:0] alpha138_0_x_locator0;
  wire [9:0] alpha138_1_x_locator1;
  wire [9:0] alpha138_2_x_locator2;
  wire [9:0] alpha138_3_x_locator3;
  wire [9:0] alpha139_0_x_locator0;
  wire [9:0] alpha139_1_x_locator1;
  wire [9:0] alpha139_2_x_locator2;
  wire [9:0] alpha139_3_x_locator3;
  wire [9:0] alpha140_0_x_locator0;
  wire [9:0] alpha140_1_x_locator1;
  wire [9:0] alpha140_2_x_locator2;
  wire [9:0] alpha140_3_x_locator3;
  wire [9:0] alpha141_0_x_locator0;
  wire [9:0] alpha141_1_x_locator1;
  wire [9:0] alpha141_2_x_locator2;
  wire [9:0] alpha141_3_x_locator3;
  wire [9:0] alpha142_0_x_locator0;
  wire [9:0] alpha142_1_x_locator1;
  wire [9:0] alpha142_2_x_locator2;
  wire [9:0] alpha142_3_x_locator3;
  wire [9:0] alpha143_0_x_locator0;
  wire [9:0] alpha143_1_x_locator1;
  wire [9:0] alpha143_2_x_locator2;
  wire [9:0] alpha143_3_x_locator3;
  wire [9:0] alpha144_0_x_locator0;
  wire [9:0] alpha144_1_x_locator1;
  wire [9:0] alpha144_2_x_locator2;
  wire [9:0] alpha144_3_x_locator3;
  wire [9:0] alpha145_0_x_locator0;
  wire [9:0] alpha145_1_x_locator1;
  wire [9:0] alpha145_2_x_locator2;
  wire [9:0] alpha145_3_x_locator3;
  wire [9:0] alpha146_0_x_locator0;
  wire [9:0] alpha146_1_x_locator1;
  wire [9:0] alpha146_2_x_locator2;
  wire [9:0] alpha146_3_x_locator3;
  wire [9:0] alpha147_0_x_locator0;
  wire [9:0] alpha147_1_x_locator1;
  wire [9:0] alpha147_2_x_locator2;
  wire [9:0] alpha147_3_x_locator3;
  wire [9:0] alpha148_0_x_locator0;
  wire [9:0] alpha148_1_x_locator1;
  wire [9:0] alpha148_2_x_locator2;
  wire [9:0] alpha148_3_x_locator3;
  wire [9:0] alpha149_0_x_locator0;
  wire [9:0] alpha149_1_x_locator1;
  wire [9:0] alpha149_2_x_locator2;
  wire [9:0] alpha149_3_x_locator3;
  wire [9:0] alpha150_0_x_locator0;
  wire [9:0] alpha150_1_x_locator1;
  wire [9:0] alpha150_2_x_locator2;
  wire [9:0] alpha150_3_x_locator3;
  wire [9:0] alpha151_0_x_locator0;
  wire [9:0] alpha151_1_x_locator1;
  wire [9:0] alpha151_2_x_locator2;
  wire [9:0] alpha151_3_x_locator3;
  wire [9:0] alpha152_0_x_locator0;
  wire [9:0] alpha152_1_x_locator1;
  wire [9:0] alpha152_2_x_locator2;
  wire [9:0] alpha152_3_x_locator3;
  wire [9:0] alpha153_0_x_locator0;
  wire [9:0] alpha153_1_x_locator1;
  wire [9:0] alpha153_2_x_locator2;
  wire [9:0] alpha153_3_x_locator3;
  wire [9:0] alpha154_0_x_locator0;
  wire [9:0] alpha154_1_x_locator1;
  wire [9:0] alpha154_2_x_locator2;
  wire [9:0] alpha154_3_x_locator3;
  wire [9:0] alpha155_0_x_locator0;
  wire [9:0] alpha155_1_x_locator1;
  wire [9:0] alpha155_2_x_locator2;
  wire [9:0] alpha155_3_x_locator3;
  wire [9:0] alpha156_0_x_locator0;
  wire [9:0] alpha156_1_x_locator1;
  wire [9:0] alpha156_2_x_locator2;
  wire [9:0] alpha156_3_x_locator3;
  wire [9:0] alpha157_0_x_locator0;
  wire [9:0] alpha157_1_x_locator1;
  wire [9:0] alpha157_2_x_locator2;
  wire [9:0] alpha157_3_x_locator3;
  wire [9:0] alpha158_0_x_locator0;
  wire [9:0] alpha158_1_x_locator1;
  wire [9:0] alpha158_2_x_locator2;
  wire [9:0] alpha158_3_x_locator3;
  wire [9:0] alpha159_0_x_locator0;
  wire [9:0] alpha159_1_x_locator1;
  wire [9:0] alpha159_2_x_locator2;
  wire [9:0] alpha159_3_x_locator3;
  wire [9:0] alpha160_0_x_locator0;
  wire [9:0] alpha160_1_x_locator1;
  wire [9:0] alpha160_2_x_locator2;
  wire [9:0] alpha160_3_x_locator3;
  wire [9:0] alpha161_0_x_locator0;
  wire [9:0] alpha161_1_x_locator1;
  wire [9:0] alpha161_2_x_locator2;
  wire [9:0] alpha161_3_x_locator3;
  wire [9:0] alpha162_0_x_locator0;
  wire [9:0] alpha162_1_x_locator1;
  wire [9:0] alpha162_2_x_locator2;
  wire [9:0] alpha162_3_x_locator3;
  wire [9:0] alpha163_0_x_locator0;
  wire [9:0] alpha163_1_x_locator1;
  wire [9:0] alpha163_2_x_locator2;
  wire [9:0] alpha163_3_x_locator3;
  wire [9:0] alpha164_0_x_locator0;
  wire [9:0] alpha164_1_x_locator1;
  wire [9:0] alpha164_2_x_locator2;
  wire [9:0] alpha164_3_x_locator3;
  wire [9:0] alpha165_0_x_locator0;
  wire [9:0] alpha165_1_x_locator1;
  wire [9:0] alpha165_2_x_locator2;
  wire [9:0] alpha165_3_x_locator3;
  wire [9:0] alpha166_0_x_locator0;
  wire [9:0] alpha166_1_x_locator1;
  wire [9:0] alpha166_2_x_locator2;
  wire [9:0] alpha166_3_x_locator3;
  wire [9:0] alpha167_0_x_locator0;
  wire [9:0] alpha167_1_x_locator1;
  wire [9:0] alpha167_2_x_locator2;
  wire [9:0] alpha167_3_x_locator3;
  wire [9:0] alpha168_0_x_locator0;
  wire [9:0] alpha168_1_x_locator1;
  wire [9:0] alpha168_2_x_locator2;
  wire [9:0] alpha168_3_x_locator3;
  wire [9:0] alpha169_0_x_locator0;
  wire [9:0] alpha169_1_x_locator1;
  wire [9:0] alpha169_2_x_locator2;
  wire [9:0] alpha169_3_x_locator3;
  wire [9:0] alpha170_0_x_locator0;
  wire [9:0] alpha170_1_x_locator1;
  wire [9:0] alpha170_2_x_locator2;
  wire [9:0] alpha170_3_x_locator3;
  wire [9:0] alpha171_0_x_locator0;
  wire [9:0] alpha171_1_x_locator1;
  wire [9:0] alpha171_2_x_locator2;
  wire [9:0] alpha171_3_x_locator3;
  wire [9:0] alpha172_0_x_locator0;
  wire [9:0] alpha172_1_x_locator1;
  wire [9:0] alpha172_2_x_locator2;
  wire [9:0] alpha172_3_x_locator3;
  wire [9:0] alpha173_0_x_locator0;
  wire [9:0] alpha173_1_x_locator1;
  wire [9:0] alpha173_2_x_locator2;
  wire [9:0] alpha173_3_x_locator3;
  wire [9:0] alpha174_0_x_locator0;
  wire [9:0] alpha174_1_x_locator1;
  wire [9:0] alpha174_2_x_locator2;
  wire [9:0] alpha174_3_x_locator3;
  wire [9:0] alpha175_0_x_locator0;
  wire [9:0] alpha175_1_x_locator1;
  wire [9:0] alpha175_2_x_locator2;
  wire [9:0] alpha175_3_x_locator3;
  wire [9:0] alpha176_0_x_locator0;
  wire [9:0] alpha176_1_x_locator1;
  wire [9:0] alpha176_2_x_locator2;
  wire [9:0] alpha176_3_x_locator3;
  wire [9:0] alpha177_0_x_locator0;
  wire [9:0] alpha177_1_x_locator1;
  wire [9:0] alpha177_2_x_locator2;
  wire [9:0] alpha177_3_x_locator3;
  wire [9:0] alpha178_0_x_locator0;
  wire [9:0] alpha178_1_x_locator1;
  wire [9:0] alpha178_2_x_locator2;
  wire [9:0] alpha178_3_x_locator3;
  wire [9:0] alpha179_0_x_locator0;
  wire [9:0] alpha179_1_x_locator1;
  wire [9:0] alpha179_2_x_locator2;
  wire [9:0] alpha179_3_x_locator3;
  wire [9:0] alpha180_0_x_locator0;
  wire [9:0] alpha180_1_x_locator1;
  wire [9:0] alpha180_2_x_locator2;
  wire [9:0] alpha180_3_x_locator3;
  wire [9:0] alpha181_0_x_locator0;
  wire [9:0] alpha181_1_x_locator1;
  wire [9:0] alpha181_2_x_locator2;
  wire [9:0] alpha181_3_x_locator3;
  wire [9:0] alpha182_0_x_locator0;
  wire [9:0] alpha182_1_x_locator1;
  wire [9:0] alpha182_2_x_locator2;
  wire [9:0] alpha182_3_x_locator3;
  wire [9:0] alpha183_0_x_locator0;
  wire [9:0] alpha183_1_x_locator1;
  wire [9:0] alpha183_2_x_locator2;
  wire [9:0] alpha183_3_x_locator3;
  wire [9:0] alpha184_0_x_locator0;
  wire [9:0] alpha184_1_x_locator1;
  wire [9:0] alpha184_2_x_locator2;
  wire [9:0] alpha184_3_x_locator3;
  wire [9:0] alpha185_0_x_locator0;
  wire [9:0] alpha185_1_x_locator1;
  wire [9:0] alpha185_2_x_locator2;
  wire [9:0] alpha185_3_x_locator3;
  wire [9:0] alpha186_0_x_locator0;
  wire [9:0] alpha186_1_x_locator1;
  wire [9:0] alpha186_2_x_locator2;
  wire [9:0] alpha186_3_x_locator3;
  wire [9:0] alpha187_0_x_locator0;
  wire [9:0] alpha187_1_x_locator1;
  wire [9:0] alpha187_2_x_locator2;
  wire [9:0] alpha187_3_x_locator3;
  wire [9:0] alpha188_0_x_locator0;
  wire [9:0] alpha188_1_x_locator1;
  wire [9:0] alpha188_2_x_locator2;
  wire [9:0] alpha188_3_x_locator3;
  wire [9:0] alpha189_0_x_locator0;
  wire [9:0] alpha189_1_x_locator1;
  wire [9:0] alpha189_2_x_locator2;
  wire [9:0] alpha189_3_x_locator3;
  wire [9:0] alpha190_0_x_locator0;
  wire [9:0] alpha190_1_x_locator1;
  wire [9:0] alpha190_2_x_locator2;
  wire [9:0] alpha190_3_x_locator3;
  wire [9:0] alpha191_0_x_locator0;
  wire [9:0] alpha191_1_x_locator1;
  wire [9:0] alpha191_2_x_locator2;
  wire [9:0] alpha191_3_x_locator3;
  wire [9:0] alpha192_0_x_locator0;
  wire [9:0] alpha192_1_x_locator1;
  wire [9:0] alpha192_2_x_locator2;
  wire [9:0] alpha192_3_x_locator3;
  wire [9:0] alpha193_0_x_locator0;
  wire [9:0] alpha193_1_x_locator1;
  wire [9:0] alpha193_2_x_locator2;
  wire [9:0] alpha193_3_x_locator3;
  wire [9:0] alpha194_0_x_locator0;
  wire [9:0] alpha194_1_x_locator1;
  wire [9:0] alpha194_2_x_locator2;
  wire [9:0] alpha194_3_x_locator3;
  wire [9:0] alpha195_0_x_locator0;
  wire [9:0] alpha195_1_x_locator1;
  wire [9:0] alpha195_2_x_locator2;
  wire [9:0] alpha195_3_x_locator3;
  wire [9:0] alpha196_0_x_locator0;
  wire [9:0] alpha196_1_x_locator1;
  wire [9:0] alpha196_2_x_locator2;
  wire [9:0] alpha196_3_x_locator3;
  wire [9:0] alpha197_0_x_locator0;
  wire [9:0] alpha197_1_x_locator1;
  wire [9:0] alpha197_2_x_locator2;
  wire [9:0] alpha197_3_x_locator3;
  wire [9:0] alpha198_0_x_locator0;
  wire [9:0] alpha198_1_x_locator1;
  wire [9:0] alpha198_2_x_locator2;
  wire [9:0] alpha198_3_x_locator3;
  wire [9:0] alpha199_0_x_locator0;
  wire [9:0] alpha199_1_x_locator1;
  wire [9:0] alpha199_2_x_locator2;
  wire [9:0] alpha199_3_x_locator3;
  wire [9:0] alpha200_0_x_locator0;
  wire [9:0] alpha200_1_x_locator1;
  wire [9:0] alpha200_2_x_locator2;
  wire [9:0] alpha200_3_x_locator3;
  wire [9:0] alpha201_0_x_locator0;
  wire [9:0] alpha201_1_x_locator1;
  wire [9:0] alpha201_2_x_locator2;
  wire [9:0] alpha201_3_x_locator3;
  wire [9:0] alpha202_0_x_locator0;
  wire [9:0] alpha202_1_x_locator1;
  wire [9:0] alpha202_2_x_locator2;
  wire [9:0] alpha202_3_x_locator3;
  wire [9:0] alpha203_0_x_locator0;
  wire [9:0] alpha203_1_x_locator1;
  wire [9:0] alpha203_2_x_locator2;
  wire [9:0] alpha203_3_x_locator3;
  wire [9:0] alpha204_0_x_locator0;
  wire [9:0] alpha204_1_x_locator1;
  wire [9:0] alpha204_2_x_locator2;
  wire [9:0] alpha204_3_x_locator3;
  wire [9:0] alpha205_0_x_locator0;
  wire [9:0] alpha205_1_x_locator1;
  wire [9:0] alpha205_2_x_locator2;
  wire [9:0] alpha205_3_x_locator3;
  wire [9:0] alpha206_0_x_locator0;
  wire [9:0] alpha206_1_x_locator1;
  wire [9:0] alpha206_2_x_locator2;
  wire [9:0] alpha206_3_x_locator3;
  wire [9:0] alpha207_0_x_locator0;
  wire [9:0] alpha207_1_x_locator1;
  wire [9:0] alpha207_2_x_locator2;
  wire [9:0] alpha207_3_x_locator3;
  wire [9:0] alpha208_0_x_locator0;
  wire [9:0] alpha208_1_x_locator1;
  wire [9:0] alpha208_2_x_locator2;
  wire [9:0] alpha208_3_x_locator3;
  wire [9:0] alpha209_0_x_locator0;
  wire [9:0] alpha209_1_x_locator1;
  wire [9:0] alpha209_2_x_locator2;
  wire [9:0] alpha209_3_x_locator3;
  wire [9:0] alpha210_0_x_locator0;
  wire [9:0] alpha210_1_x_locator1;
  wire [9:0] alpha210_2_x_locator2;
  wire [9:0] alpha210_3_x_locator3;
  wire [9:0] alpha211_0_x_locator0;
  wire [9:0] alpha211_1_x_locator1;
  wire [9:0] alpha211_2_x_locator2;
  wire [9:0] alpha211_3_x_locator3;
  wire [9:0] alpha212_0_x_locator0;
  wire [9:0] alpha212_1_x_locator1;
  wire [9:0] alpha212_2_x_locator2;
  wire [9:0] alpha212_3_x_locator3;
  wire [9:0] alpha213_0_x_locator0;
  wire [9:0] alpha213_1_x_locator1;
  wire [9:0] alpha213_2_x_locator2;
  wire [9:0] alpha213_3_x_locator3;
  wire [9:0] alpha214_0_x_locator0;
  wire [9:0] alpha214_1_x_locator1;
  wire [9:0] alpha214_2_x_locator2;
  wire [9:0] alpha214_3_x_locator3;
  wire [9:0] alpha215_0_x_locator0;
  wire [9:0] alpha215_1_x_locator1;
  wire [9:0] alpha215_2_x_locator2;
  wire [9:0] alpha215_3_x_locator3;
  wire [9:0] alpha216_0_x_locator0;
  wire [9:0] alpha216_1_x_locator1;
  wire [9:0] alpha216_2_x_locator2;
  wire [9:0] alpha216_3_x_locator3;
  wire [9:0] alpha217_0_x_locator0;
  wire [9:0] alpha217_1_x_locator1;
  wire [9:0] alpha217_2_x_locator2;
  wire [9:0] alpha217_3_x_locator3;
  wire [9:0] alpha218_0_x_locator0;
  wire [9:0] alpha218_1_x_locator1;
  wire [9:0] alpha218_2_x_locator2;
  wire [9:0] alpha218_3_x_locator3;
  wire [9:0] alpha219_0_x_locator0;
  wire [9:0] alpha219_1_x_locator1;
  wire [9:0] alpha219_2_x_locator2;
  wire [9:0] alpha219_3_x_locator3;
  wire [9:0] alpha220_0_x_locator0;
  wire [9:0] alpha220_1_x_locator1;
  wire [9:0] alpha220_2_x_locator2;
  wire [9:0] alpha220_3_x_locator3;
  wire [9:0] alpha221_0_x_locator0;
  wire [9:0] alpha221_1_x_locator1;
  wire [9:0] alpha221_2_x_locator2;
  wire [9:0] alpha221_3_x_locator3;
  wire [9:0] alpha222_0_x_locator0;
  wire [9:0] alpha222_1_x_locator1;
  wire [9:0] alpha222_2_x_locator2;
  wire [9:0] alpha222_3_x_locator3;
  wire [9:0] alpha223_0_x_locator0;
  wire [9:0] alpha223_1_x_locator1;
  wire [9:0] alpha223_2_x_locator2;
  wire [9:0] alpha223_3_x_locator3;
  wire [9:0] alpha224_0_x_locator0;
  wire [9:0] alpha224_1_x_locator1;
  wire [9:0] alpha224_2_x_locator2;
  wire [9:0] alpha224_3_x_locator3;
  wire [9:0] alpha225_0_x_locator0;
  wire [9:0] alpha225_1_x_locator1;
  wire [9:0] alpha225_2_x_locator2;
  wire [9:0] alpha225_3_x_locator3;
  wire [9:0] alpha226_0_x_locator0;
  wire [9:0] alpha226_1_x_locator1;
  wire [9:0] alpha226_2_x_locator2;
  wire [9:0] alpha226_3_x_locator3;
  wire [9:0] alpha227_0_x_locator0;
  wire [9:0] alpha227_1_x_locator1;
  wire [9:0] alpha227_2_x_locator2;
  wire [9:0] alpha227_3_x_locator3;
  wire [9:0] alpha228_0_x_locator0;
  wire [9:0] alpha228_1_x_locator1;
  wire [9:0] alpha228_2_x_locator2;
  wire [9:0] alpha228_3_x_locator3;
  wire [9:0] alpha229_0_x_locator0;
  wire [9:0] alpha229_1_x_locator1;
  wire [9:0] alpha229_2_x_locator2;
  wire [9:0] alpha229_3_x_locator3;
  wire [9:0] alpha230_0_x_locator0;
  wire [9:0] alpha230_1_x_locator1;
  wire [9:0] alpha230_2_x_locator2;
  wire [9:0] alpha230_3_x_locator3;
  wire [9:0] alpha231_0_x_locator0;
  wire [9:0] alpha231_1_x_locator1;
  wire [9:0] alpha231_2_x_locator2;
  wire [9:0] alpha231_3_x_locator3;
  wire [9:0] alpha232_0_x_locator0;
  wire [9:0] alpha232_1_x_locator1;
  wire [9:0] alpha232_2_x_locator2;
  wire [9:0] alpha232_3_x_locator3;
  wire [9:0] alpha233_0_x_locator0;
  wire [9:0] alpha233_1_x_locator1;
  wire [9:0] alpha233_2_x_locator2;
  wire [9:0] alpha233_3_x_locator3;
  wire [9:0] alpha234_0_x_locator0;
  wire [9:0] alpha234_1_x_locator1;
  wire [9:0] alpha234_2_x_locator2;
  wire [9:0] alpha234_3_x_locator3;
  wire [9:0] alpha235_0_x_locator0;
  wire [9:0] alpha235_1_x_locator1;
  wire [9:0] alpha235_2_x_locator2;
  wire [9:0] alpha235_3_x_locator3;
  wire [9:0] alpha236_0_x_locator0;
  wire [9:0] alpha236_1_x_locator1;
  wire [9:0] alpha236_2_x_locator2;
  wire [9:0] alpha236_3_x_locator3;
  wire [9:0] alpha237_0_x_locator0;
  wire [9:0] alpha237_1_x_locator1;
  wire [9:0] alpha237_2_x_locator2;
  wire [9:0] alpha237_3_x_locator3;
  wire [9:0] alpha238_0_x_locator0;
  wire [9:0] alpha238_1_x_locator1;
  wire [9:0] alpha238_2_x_locator2;
  wire [9:0] alpha238_3_x_locator3;
  wire [9:0] alpha239_0_x_locator0;
  wire [9:0] alpha239_1_x_locator1;
  wire [9:0] alpha239_2_x_locator2;
  wire [9:0] alpha239_3_x_locator3;
  wire [9:0] alpha240_0_x_locator0;
  wire [9:0] alpha240_1_x_locator1;
  wire [9:0] alpha240_2_x_locator2;
  wire [9:0] alpha240_3_x_locator3;
  wire [9:0] alpha241_0_x_locator0;
  wire [9:0] alpha241_1_x_locator1;
  wire [9:0] alpha241_2_x_locator2;
  wire [9:0] alpha241_3_x_locator3;
  wire [9:0] alpha242_0_x_locator0;
  wire [9:0] alpha242_1_x_locator1;
  wire [9:0] alpha242_2_x_locator2;
  wire [9:0] alpha242_3_x_locator3;
  wire [9:0] alpha243_0_x_locator0;
  wire [9:0] alpha243_1_x_locator1;
  wire [9:0] alpha243_2_x_locator2;
  wire [9:0] alpha243_3_x_locator3;
  wire [9:0] alpha244_0_x_locator0;
  wire [9:0] alpha244_1_x_locator1;
  wire [9:0] alpha244_2_x_locator2;
  wire [9:0] alpha244_3_x_locator3;
  wire [9:0] alpha245_0_x_locator0;
  wire [9:0] alpha245_1_x_locator1;
  wire [9:0] alpha245_2_x_locator2;
  wire [9:0] alpha245_3_x_locator3;
  wire [9:0] alpha246_0_x_locator0;
  wire [9:0] alpha246_1_x_locator1;
  wire [9:0] alpha246_2_x_locator2;
  wire [9:0] alpha246_3_x_locator3;
  wire [9:0] alpha247_0_x_locator0;
  wire [9:0] alpha247_1_x_locator1;
  wire [9:0] alpha247_2_x_locator2;
  wire [9:0] alpha247_3_x_locator3;
  wire [9:0] alpha248_0_x_locator0;
  wire [9:0] alpha248_1_x_locator1;
  wire [9:0] alpha248_2_x_locator2;
  wire [9:0] alpha248_3_x_locator3;
  wire [9:0] alpha249_0_x_locator0;
  wire [9:0] alpha249_1_x_locator1;
  wire [9:0] alpha249_2_x_locator2;
  wire [9:0] alpha249_3_x_locator3;
  wire [9:0] alpha250_0_x_locator0;
  wire [9:0] alpha250_1_x_locator1;
  wire [9:0] alpha250_2_x_locator2;
  wire [9:0] alpha250_3_x_locator3;
  wire [9:0] alpha251_0_x_locator0;
  wire [9:0] alpha251_1_x_locator1;
  wire [9:0] alpha251_2_x_locator2;
  wire [9:0] alpha251_3_x_locator3;
  wire [9:0] alpha252_0_x_locator0;
  wire [9:0] alpha252_1_x_locator1;
  wire [9:0] alpha252_2_x_locator2;
  wire [9:0] alpha252_3_x_locator3;
  wire [9:0] alpha253_0_x_locator0;
  wire [9:0] alpha253_1_x_locator1;
  wire [9:0] alpha253_2_x_locator2;
  wire [9:0] alpha253_3_x_locator3;
  wire [9:0] alpha254_0_x_locator0;
  wire [9:0] alpha254_1_x_locator1;
  wire [9:0] alpha254_2_x_locator2;
  wire [9:0] alpha254_3_x_locator3;
  wire [9:0] alpha255_0_x_locator0;
  wire [9:0] alpha255_1_x_locator1;
  wire [9:0] alpha255_2_x_locator2;
  wire [9:0] alpha255_3_x_locator3;
  wire [9:0] alpha256_0_x_locator0;
  wire [9:0] alpha256_1_x_locator1;
  wire [9:0] alpha256_2_x_locator2;
  wire [9:0] alpha256_3_x_locator3;
  wire [9:0] alpha257_0_x_locator0;
  wire [9:0] alpha257_1_x_locator1;
  wire [9:0] alpha257_2_x_locator2;
  wire [9:0] alpha257_3_x_locator3;
  wire [9:0] alpha258_0_x_locator0;
  wire [9:0] alpha258_1_x_locator1;
  wire [9:0] alpha258_2_x_locator2;
  wire [9:0] alpha258_3_x_locator3;
  wire [9:0] alpha259_0_x_locator0;
  wire [9:0] alpha259_1_x_locator1;
  wire [9:0] alpha259_2_x_locator2;
  wire [9:0] alpha259_3_x_locator3;
  wire [9:0] alpha260_0_x_locator0;
  wire [9:0] alpha260_1_x_locator1;
  wire [9:0] alpha260_2_x_locator2;
  wire [9:0] alpha260_3_x_locator3;
  wire [9:0] alpha261_0_x_locator0;
  wire [9:0] alpha261_1_x_locator1;
  wire [9:0] alpha261_2_x_locator2;
  wire [9:0] alpha261_3_x_locator3;
  wire [9:0] alpha262_0_x_locator0;
  wire [9:0] alpha262_1_x_locator1;
  wire [9:0] alpha262_2_x_locator2;
  wire [9:0] alpha262_3_x_locator3;
  wire [9:0] alpha263_0_x_locator0;
  wire [9:0] alpha263_1_x_locator1;
  wire [9:0] alpha263_2_x_locator2;
  wire [9:0] alpha263_3_x_locator3;
  wire [9:0] alpha264_0_x_locator0;
  wire [9:0] alpha264_1_x_locator1;
  wire [9:0] alpha264_2_x_locator2;
  wire [9:0] alpha264_3_x_locator3;
  wire [9:0] alpha265_0_x_locator0;
  wire [9:0] alpha265_1_x_locator1;
  wire [9:0] alpha265_2_x_locator2;
  wire [9:0] alpha265_3_x_locator3;
  wire [9:0] alpha266_0_x_locator0;
  wire [9:0] alpha266_1_x_locator1;
  wire [9:0] alpha266_2_x_locator2;
  wire [9:0] alpha266_3_x_locator3;
  wire [9:0] alpha267_0_x_locator0;
  wire [9:0] alpha267_1_x_locator1;
  wire [9:0] alpha267_2_x_locator2;
  wire [9:0] alpha267_3_x_locator3;
  wire [9:0] alpha268_0_x_locator0;
  wire [9:0] alpha268_1_x_locator1;
  wire [9:0] alpha268_2_x_locator2;
  wire [9:0] alpha268_3_x_locator3;
  wire [9:0] alpha269_0_x_locator0;
  wire [9:0] alpha269_1_x_locator1;
  wire [9:0] alpha269_2_x_locator2;
  wire [9:0] alpha269_3_x_locator3;
  wire [9:0] alpha270_0_x_locator0;
  wire [9:0] alpha270_1_x_locator1;
  wire [9:0] alpha270_2_x_locator2;
  wire [9:0] alpha270_3_x_locator3;
  wire [9:0] alpha271_0_x_locator0;
  wire [9:0] alpha271_1_x_locator1;
  wire [9:0] alpha271_2_x_locator2;
  wire [9:0] alpha271_3_x_locator3;
  wire [9:0] alpha272_0_x_locator0;
  wire [9:0] alpha272_1_x_locator1;
  wire [9:0] alpha272_2_x_locator2;
  wire [9:0] alpha272_3_x_locator3;
  wire [9:0] alpha273_0_x_locator0;
  wire [9:0] alpha273_1_x_locator1;
  wire [9:0] alpha273_2_x_locator2;
  wire [9:0] alpha273_3_x_locator3;
  wire [9:0] alpha274_0_x_locator0;
  wire [9:0] alpha274_1_x_locator1;
  wire [9:0] alpha274_2_x_locator2;
  wire [9:0] alpha274_3_x_locator3;
  wire [9:0] alpha275_0_x_locator0;
  wire [9:0] alpha275_1_x_locator1;
  wire [9:0] alpha275_2_x_locator2;
  wire [9:0] alpha275_3_x_locator3;
  wire [9:0] alpha276_0_x_locator0;
  wire [9:0] alpha276_1_x_locator1;
  wire [9:0] alpha276_2_x_locator2;
  wire [9:0] alpha276_3_x_locator3;
  wire [9:0] alpha277_0_x_locator0;
  wire [9:0] alpha277_1_x_locator1;
  wire [9:0] alpha277_2_x_locator2;
  wire [9:0] alpha277_3_x_locator3;
  wire [9:0] alpha278_0_x_locator0;
  wire [9:0] alpha278_1_x_locator1;
  wire [9:0] alpha278_2_x_locator2;
  wire [9:0] alpha278_3_x_locator3;
  wire [9:0] alpha279_0_x_locator0;
  wire [9:0] alpha279_1_x_locator1;
  wire [9:0] alpha279_2_x_locator2;
  wire [9:0] alpha279_3_x_locator3;
  wire [9:0] alpha280_0_x_locator0;
  wire [9:0] alpha280_1_x_locator1;
  wire [9:0] alpha280_2_x_locator2;
  wire [9:0] alpha280_3_x_locator3;
  wire [9:0] alpha281_0_x_locator0;
  wire [9:0] alpha281_1_x_locator1;
  wire [9:0] alpha281_2_x_locator2;
  wire [9:0] alpha281_3_x_locator3;
  wire [9:0] alpha282_0_x_locator0;
  wire [9:0] alpha282_1_x_locator1;
  wire [9:0] alpha282_2_x_locator2;
  wire [9:0] alpha282_3_x_locator3;
  wire [9:0] alpha283_0_x_locator0;
  wire [9:0] alpha283_1_x_locator1;
  wire [9:0] alpha283_2_x_locator2;
  wire [9:0] alpha283_3_x_locator3;
  wire [9:0] alpha284_0_x_locator0;
  wire [9:0] alpha284_1_x_locator1;
  wire [9:0] alpha284_2_x_locator2;
  wire [9:0] alpha284_3_x_locator3;
  wire [9:0] alpha285_0_x_locator0;
  wire [9:0] alpha285_1_x_locator1;
  wire [9:0] alpha285_2_x_locator2;
  wire [9:0] alpha285_3_x_locator3;
  wire [9:0] alpha286_0_x_locator0;
  wire [9:0] alpha286_1_x_locator1;
  wire [9:0] alpha286_2_x_locator2;
  wire [9:0] alpha286_3_x_locator3;
  wire [9:0] alpha287_0_x_locator0;
  wire [9:0] alpha287_1_x_locator1;
  wire [9:0] alpha287_2_x_locator2;
  wire [9:0] alpha287_3_x_locator3;
  wire [9:0] alpha288_0_x_locator0;
  wire [9:0] alpha288_1_x_locator1;
  wire [9:0] alpha288_2_x_locator2;
  wire [9:0] alpha288_3_x_locator3;
  wire [9:0] alpha289_0_x_locator0;
  wire [9:0] alpha289_1_x_locator1;
  wire [9:0] alpha289_2_x_locator2;
  wire [9:0] alpha289_3_x_locator3;
  wire [9:0] alpha290_0_x_locator0;
  wire [9:0] alpha290_1_x_locator1;
  wire [9:0] alpha290_2_x_locator2;
  wire [9:0] alpha290_3_x_locator3;
  wire [9:0] alpha291_0_x_locator0;
  wire [9:0] alpha291_1_x_locator1;
  wire [9:0] alpha291_2_x_locator2;
  wire [9:0] alpha291_3_x_locator3;
  wire [9:0] alpha292_0_x_locator0;
  wire [9:0] alpha292_1_x_locator1;
  wire [9:0] alpha292_2_x_locator2;
  wire [9:0] alpha292_3_x_locator3;
  wire [9:0] alpha293_0_x_locator0;
  wire [9:0] alpha293_1_x_locator1;
  wire [9:0] alpha293_2_x_locator2;
  wire [9:0] alpha293_3_x_locator3;
  wire [9:0] alpha294_0_x_locator0;
  wire [9:0] alpha294_1_x_locator1;
  wire [9:0] alpha294_2_x_locator2;
  wire [9:0] alpha294_3_x_locator3;
  wire [9:0] alpha295_0_x_locator0;
  wire [9:0] alpha295_1_x_locator1;
  wire [9:0] alpha295_2_x_locator2;
  wire [9:0] alpha295_3_x_locator3;
  wire [9:0] alpha296_0_x_locator0;
  wire [9:0] alpha296_1_x_locator1;
  wire [9:0] alpha296_2_x_locator2;
  wire [9:0] alpha296_3_x_locator3;
  wire [9:0] alpha297_0_x_locator0;
  wire [9:0] alpha297_1_x_locator1;
  wire [9:0] alpha297_2_x_locator2;
  wire [9:0] alpha297_3_x_locator3;
  wire [9:0] alpha298_0_x_locator0;
  wire [9:0] alpha298_1_x_locator1;
  wire [9:0] alpha298_2_x_locator2;
  wire [9:0] alpha298_3_x_locator3;
  wire [9:0] alpha299_0_x_locator0;
  wire [9:0] alpha299_1_x_locator1;
  wire [9:0] alpha299_2_x_locator2;
  wire [9:0] alpha299_3_x_locator3;
  wire [9:0] alpha300_0_x_locator0;
  wire [9:0] alpha300_1_x_locator1;
  wire [9:0] alpha300_2_x_locator2;
  wire [9:0] alpha300_3_x_locator3;
  wire [9:0] alpha301_0_x_locator0;
  wire [9:0] alpha301_1_x_locator1;
  wire [9:0] alpha301_2_x_locator2;
  wire [9:0] alpha301_3_x_locator3;
  wire [9:0] alpha302_0_x_locator0;
  wire [9:0] alpha302_1_x_locator1;
  wire [9:0] alpha302_2_x_locator2;
  wire [9:0] alpha302_3_x_locator3;
  wire [9:0] alpha303_0_x_locator0;
  wire [9:0] alpha303_1_x_locator1;
  wire [9:0] alpha303_2_x_locator2;
  wire [9:0] alpha303_3_x_locator3;
  wire [9:0] alpha304_0_x_locator0;
  wire [9:0] alpha304_1_x_locator1;
  wire [9:0] alpha304_2_x_locator2;
  wire [9:0] alpha304_3_x_locator3;
  wire [9:0] alpha305_0_x_locator0;
  wire [9:0] alpha305_1_x_locator1;
  wire [9:0] alpha305_2_x_locator2;
  wire [9:0] alpha305_3_x_locator3;
  wire [9:0] alpha306_0_x_locator0;
  wire [9:0] alpha306_1_x_locator1;
  wire [9:0] alpha306_2_x_locator2;
  wire [9:0] alpha306_3_x_locator3;
  wire [9:0] alpha307_0_x_locator0;
  wire [9:0] alpha307_1_x_locator1;
  wire [9:0] alpha307_2_x_locator2;
  wire [9:0] alpha307_3_x_locator3;
  wire [9:0] alpha308_0_x_locator0;
  wire [9:0] alpha308_1_x_locator1;
  wire [9:0] alpha308_2_x_locator2;
  wire [9:0] alpha308_3_x_locator3;
  wire [9:0] alpha309_0_x_locator0;
  wire [9:0] alpha309_1_x_locator1;
  wire [9:0] alpha309_2_x_locator2;
  wire [9:0] alpha309_3_x_locator3;
  wire [9:0] alpha310_0_x_locator0;
  wire [9:0] alpha310_1_x_locator1;
  wire [9:0] alpha310_2_x_locator2;
  wire [9:0] alpha310_3_x_locator3;
  wire [9:0] alpha311_0_x_locator0;
  wire [9:0] alpha311_1_x_locator1;
  wire [9:0] alpha311_2_x_locator2;
  wire [9:0] alpha311_3_x_locator3;
  wire [9:0] alpha312_0_x_locator0;
  wire [9:0] alpha312_1_x_locator1;
  wire [9:0] alpha312_2_x_locator2;
  wire [9:0] alpha312_3_x_locator3;
  wire [9:0] alpha313_0_x_locator0;
  wire [9:0] alpha313_1_x_locator1;
  wire [9:0] alpha313_2_x_locator2;
  wire [9:0] alpha313_3_x_locator3;
  wire [9:0] alpha314_0_x_locator0;
  wire [9:0] alpha314_1_x_locator1;
  wire [9:0] alpha314_2_x_locator2;
  wire [9:0] alpha314_3_x_locator3;
  wire [9:0] alpha315_0_x_locator0;
  wire [9:0] alpha315_1_x_locator1;
  wire [9:0] alpha315_2_x_locator2;
  wire [9:0] alpha315_3_x_locator3;
  wire [9:0] alpha316_0_x_locator0;
  wire [9:0] alpha316_1_x_locator1;
  wire [9:0] alpha316_2_x_locator2;
  wire [9:0] alpha316_3_x_locator3;
  wire [9:0] alpha317_0_x_locator0;
  wire [9:0] alpha317_1_x_locator1;
  wire [9:0] alpha317_2_x_locator2;
  wire [9:0] alpha317_3_x_locator3;
  wire [9:0] alpha318_0_x_locator0;
  wire [9:0] alpha318_1_x_locator1;
  wire [9:0] alpha318_2_x_locator2;
  wire [9:0] alpha318_3_x_locator3;
  wire [9:0] alpha319_0_x_locator0;
  wire [9:0] alpha319_1_x_locator1;
  wire [9:0] alpha319_2_x_locator2;
  wire [9:0] alpha319_3_x_locator3;
  wire [9:0] alpha320_0_x_locator0;
  wire [9:0] alpha320_1_x_locator1;
  wire [9:0] alpha320_2_x_locator2;
  wire [9:0] alpha320_3_x_locator3;
  wire [9:0] alpha321_0_x_locator0;
  wire [9:0] alpha321_1_x_locator1;
  wire [9:0] alpha321_2_x_locator2;
  wire [9:0] alpha321_3_x_locator3;
  wire [9:0] alpha322_0_x_locator0;
  wire [9:0] alpha322_1_x_locator1;
  wire [9:0] alpha322_2_x_locator2;
  wire [9:0] alpha322_3_x_locator3;
  wire [9:0] alpha323_0_x_locator0;
  wire [9:0] alpha323_1_x_locator1;
  wire [9:0] alpha323_2_x_locator2;
  wire [9:0] alpha323_3_x_locator3;
  wire [9:0] alpha324_0_x_locator0;
  wire [9:0] alpha324_1_x_locator1;
  wire [9:0] alpha324_2_x_locator2;
  wire [9:0] alpha324_3_x_locator3;
  wire [9:0] alpha325_0_x_locator0;
  wire [9:0] alpha325_1_x_locator1;
  wire [9:0] alpha325_2_x_locator2;
  wire [9:0] alpha325_3_x_locator3;
  wire [9:0] alpha326_0_x_locator0;
  wire [9:0] alpha326_1_x_locator1;
  wire [9:0] alpha326_2_x_locator2;
  wire [9:0] alpha326_3_x_locator3;
  wire [9:0] alpha327_0_x_locator0;
  wire [9:0] alpha327_1_x_locator1;
  wire [9:0] alpha327_2_x_locator2;
  wire [9:0] alpha327_3_x_locator3;
  wire [9:0] alpha328_0_x_locator0;
  wire [9:0] alpha328_1_x_locator1;
  wire [9:0] alpha328_2_x_locator2;
  wire [9:0] alpha328_3_x_locator3;
  wire [9:0] alpha329_0_x_locator0;
  wire [9:0] alpha329_1_x_locator1;
  wire [9:0] alpha329_2_x_locator2;
  wire [9:0] alpha329_3_x_locator3;
  wire [9:0] alpha330_0_x_locator0;
  wire [9:0] alpha330_1_x_locator1;
  wire [9:0] alpha330_2_x_locator2;
  wire [9:0] alpha330_3_x_locator3;
  wire [9:0] alpha331_0_x_locator0;
  wire [9:0] alpha331_1_x_locator1;
  wire [9:0] alpha331_2_x_locator2;
  wire [9:0] alpha331_3_x_locator3;
  wire [9:0] alpha332_0_x_locator0;
  wire [9:0] alpha332_1_x_locator1;
  wire [9:0] alpha332_2_x_locator2;
  wire [9:0] alpha332_3_x_locator3;
  wire [9:0] alpha333_0_x_locator0;
  wire [9:0] alpha333_1_x_locator1;
  wire [9:0] alpha333_2_x_locator2;
  wire [9:0] alpha333_3_x_locator3;
  wire [9:0] alpha334_0_x_locator0;
  wire [9:0] alpha334_1_x_locator1;
  wire [9:0] alpha334_2_x_locator2;
  wire [9:0] alpha334_3_x_locator3;
  wire [9:0] alpha335_0_x_locator0;
  wire [9:0] alpha335_1_x_locator1;
  wire [9:0] alpha335_2_x_locator2;
  wire [9:0] alpha335_3_x_locator3;
  wire [9:0] alpha336_0_x_locator0;
  wire [9:0] alpha336_1_x_locator1;
  wire [9:0] alpha336_2_x_locator2;
  wire [9:0] alpha336_3_x_locator3;
  wire [9:0] alpha337_0_x_locator0;
  wire [9:0] alpha337_1_x_locator1;
  wire [9:0] alpha337_2_x_locator2;
  wire [9:0] alpha337_3_x_locator3;
  wire [9:0] alpha338_0_x_locator0;
  wire [9:0] alpha338_1_x_locator1;
  wire [9:0] alpha338_2_x_locator2;
  wire [9:0] alpha338_3_x_locator3;
  wire [9:0] alpha339_0_x_locator0;
  wire [9:0] alpha339_1_x_locator1;
  wire [9:0] alpha339_2_x_locator2;
  wire [9:0] alpha339_3_x_locator3;
  wire [9:0] alpha340_0_x_locator0;
  wire [9:0] alpha340_1_x_locator1;
  wire [9:0] alpha340_2_x_locator2;
  wire [9:0] alpha340_3_x_locator3;
  wire [9:0] alpha341_0_x_locator0;
  wire [9:0] alpha341_1_x_locator1;
  wire [9:0] alpha341_2_x_locator2;
  wire [9:0] alpha341_3_x_locator3;
  wire [9:0] alpha342_0_x_locator0;
  wire [9:0] alpha342_1_x_locator1;
  wire [9:0] alpha342_2_x_locator2;
  wire [9:0] alpha342_3_x_locator3;
  wire [9:0] alpha343_0_x_locator0;
  wire [9:0] alpha343_1_x_locator1;
  wire [9:0] alpha343_2_x_locator2;
  wire [9:0] alpha343_3_x_locator3;
  wire [9:0] alpha344_0_x_locator0;
  wire [9:0] alpha344_1_x_locator1;
  wire [9:0] alpha344_2_x_locator2;
  wire [9:0] alpha344_3_x_locator3;
  wire [9:0] alpha345_0_x_locator0;
  wire [9:0] alpha345_1_x_locator1;
  wire [9:0] alpha345_2_x_locator2;
  wire [9:0] alpha345_3_x_locator3;
  wire [9:0] alpha346_0_x_locator0;
  wire [9:0] alpha346_1_x_locator1;
  wire [9:0] alpha346_2_x_locator2;
  wire [9:0] alpha346_3_x_locator3;
  wire [9:0] alpha347_0_x_locator0;
  wire [9:0] alpha347_1_x_locator1;
  wire [9:0] alpha347_2_x_locator2;
  wire [9:0] alpha347_3_x_locator3;
  wire [9:0] alpha348_0_x_locator0;
  wire [9:0] alpha348_1_x_locator1;
  wire [9:0] alpha348_2_x_locator2;
  wire [9:0] alpha348_3_x_locator3;
  wire [9:0] alpha349_0_x_locator0;
  wire [9:0] alpha349_1_x_locator1;
  wire [9:0] alpha349_2_x_locator2;
  wire [9:0] alpha349_3_x_locator3;
  wire [9:0] alpha350_0_x_locator0;
  wire [9:0] alpha350_1_x_locator1;
  wire [9:0] alpha350_2_x_locator2;
  wire [9:0] alpha350_3_x_locator3;
  wire [9:0] alpha351_0_x_locator0;
  wire [9:0] alpha351_1_x_locator1;
  wire [9:0] alpha351_2_x_locator2;
  wire [9:0] alpha351_3_x_locator3;
  wire [9:0] alpha352_0_x_locator0;
  wire [9:0] alpha352_1_x_locator1;
  wire [9:0] alpha352_2_x_locator2;
  wire [9:0] alpha352_3_x_locator3;
  wire [9:0] alpha353_0_x_locator0;
  wire [9:0] alpha353_1_x_locator1;
  wire [9:0] alpha353_2_x_locator2;
  wire [9:0] alpha353_3_x_locator3;
  wire [9:0] alpha354_0_x_locator0;
  wire [9:0] alpha354_1_x_locator1;
  wire [9:0] alpha354_2_x_locator2;
  wire [9:0] alpha354_3_x_locator3;
  wire [9:0] alpha355_0_x_locator0;
  wire [9:0] alpha355_1_x_locator1;
  wire [9:0] alpha355_2_x_locator2;
  wire [9:0] alpha355_3_x_locator3;
  wire [9:0] alpha356_0_x_locator0;
  wire [9:0] alpha356_1_x_locator1;
  wire [9:0] alpha356_2_x_locator2;
  wire [9:0] alpha356_3_x_locator3;
  wire [9:0] alpha357_0_x_locator0;
  wire [9:0] alpha357_1_x_locator1;
  wire [9:0] alpha357_2_x_locator2;
  wire [9:0] alpha357_3_x_locator3;
  wire [9:0] alpha358_0_x_locator0;
  wire [9:0] alpha358_1_x_locator1;
  wire [9:0] alpha358_2_x_locator2;
  wire [9:0] alpha358_3_x_locator3;
  wire [9:0] alpha359_0_x_locator0;
  wire [9:0] alpha359_1_x_locator1;
  wire [9:0] alpha359_2_x_locator2;
  wire [9:0] alpha359_3_x_locator3;
  wire [9:0] alpha360_0_x_locator0;
  wire [9:0] alpha360_1_x_locator1;
  wire [9:0] alpha360_2_x_locator2;
  wire [9:0] alpha360_3_x_locator3;
  wire [9:0] alpha361_0_x_locator0;
  wire [9:0] alpha361_1_x_locator1;
  wire [9:0] alpha361_2_x_locator2;
  wire [9:0] alpha361_3_x_locator3;
  wire [9:0] alpha362_0_x_locator0;
  wire [9:0] alpha362_1_x_locator1;
  wire [9:0] alpha362_2_x_locator2;
  wire [9:0] alpha362_3_x_locator3;
  wire [9:0] alpha363_0_x_locator0;
  wire [9:0] alpha363_1_x_locator1;
  wire [9:0] alpha363_2_x_locator2;
  wire [9:0] alpha363_3_x_locator3;
  wire [9:0] alpha364_0_x_locator0;
  wire [9:0] alpha364_1_x_locator1;
  wire [9:0] alpha364_2_x_locator2;
  wire [9:0] alpha364_3_x_locator3;
  wire [9:0] alpha365_0_x_locator0;
  wire [9:0] alpha365_1_x_locator1;
  wire [9:0] alpha365_2_x_locator2;
  wire [9:0] alpha365_3_x_locator3;
  wire [9:0] alpha366_0_x_locator0;
  wire [9:0] alpha366_1_x_locator1;
  wire [9:0] alpha366_2_x_locator2;
  wire [9:0] alpha366_3_x_locator3;
  wire [9:0] alpha367_0_x_locator0;
  wire [9:0] alpha367_1_x_locator1;
  wire [9:0] alpha367_2_x_locator2;
  wire [9:0] alpha367_3_x_locator3;
  wire [9:0] alpha368_0_x_locator0;
  wire [9:0] alpha368_1_x_locator1;
  wire [9:0] alpha368_2_x_locator2;
  wire [9:0] alpha368_3_x_locator3;
  wire [9:0] alpha369_0_x_locator0;
  wire [9:0] alpha369_1_x_locator1;
  wire [9:0] alpha369_2_x_locator2;
  wire [9:0] alpha369_3_x_locator3;
  wire [9:0] alpha370_0_x_locator0;
  wire [9:0] alpha370_1_x_locator1;
  wire [9:0] alpha370_2_x_locator2;
  wire [9:0] alpha370_3_x_locator3;
  wire [9:0] alpha371_0_x_locator0;
  wire [9:0] alpha371_1_x_locator1;
  wire [9:0] alpha371_2_x_locator2;
  wire [9:0] alpha371_3_x_locator3;
  wire [9:0] alpha372_0_x_locator0;
  wire [9:0] alpha372_1_x_locator1;
  wire [9:0] alpha372_2_x_locator2;
  wire [9:0] alpha372_3_x_locator3;
  wire [9:0] alpha373_0_x_locator0;
  wire [9:0] alpha373_1_x_locator1;
  wire [9:0] alpha373_2_x_locator2;
  wire [9:0] alpha373_3_x_locator3;
  wire [9:0] alpha374_0_x_locator0;
  wire [9:0] alpha374_1_x_locator1;
  wire [9:0] alpha374_2_x_locator2;
  wire [9:0] alpha374_3_x_locator3;
  wire [9:0] alpha375_0_x_locator0;
  wire [9:0] alpha375_1_x_locator1;
  wire [9:0] alpha375_2_x_locator2;
  wire [9:0] alpha375_3_x_locator3;
  wire [9:0] alpha376_0_x_locator0;
  wire [9:0] alpha376_1_x_locator1;
  wire [9:0] alpha376_2_x_locator2;
  wire [9:0] alpha376_3_x_locator3;
  wire [9:0] alpha377_0_x_locator0;
  wire [9:0] alpha377_1_x_locator1;
  wire [9:0] alpha377_2_x_locator2;
  wire [9:0] alpha377_3_x_locator3;
  wire [9:0] alpha378_0_x_locator0;
  wire [9:0] alpha378_1_x_locator1;
  wire [9:0] alpha378_2_x_locator2;
  wire [9:0] alpha378_3_x_locator3;
  wire [9:0] alpha379_0_x_locator0;
  wire [9:0] alpha379_1_x_locator1;
  wire [9:0] alpha379_2_x_locator2;
  wire [9:0] alpha379_3_x_locator3;
  wire [9:0] alpha380_0_x_locator0;
  wire [9:0] alpha380_1_x_locator1;
  wire [9:0] alpha380_2_x_locator2;
  wire [9:0] alpha380_3_x_locator3;
  wire [9:0] alpha381_0_x_locator0;
  wire [9:0] alpha381_1_x_locator1;
  wire [9:0] alpha381_2_x_locator2;
  wire [9:0] alpha381_3_x_locator3;
  wire [9:0] alpha382_0_x_locator0;
  wire [9:0] alpha382_1_x_locator1;
  wire [9:0] alpha382_2_x_locator2;
  wire [9:0] alpha382_3_x_locator3;
  wire [9:0] alpha383_0_x_locator0;
  wire [9:0] alpha383_1_x_locator1;
  wire [9:0] alpha383_2_x_locator2;
  wire [9:0] alpha383_3_x_locator3;
  wire [9:0] alpha384_0_x_locator0;
  wire [9:0] alpha384_1_x_locator1;
  wire [9:0] alpha384_2_x_locator2;
  wire [9:0] alpha384_3_x_locator3;
  wire [9:0] alpha385_0_x_locator0;
  wire [9:0] alpha385_1_x_locator1;
  wire [9:0] alpha385_2_x_locator2;
  wire [9:0] alpha385_3_x_locator3;
  wire [9:0] alpha386_0_x_locator0;
  wire [9:0] alpha386_1_x_locator1;
  wire [9:0] alpha386_2_x_locator2;
  wire [9:0] alpha386_3_x_locator3;
  wire [9:0] alpha387_0_x_locator0;
  wire [9:0] alpha387_1_x_locator1;
  wire [9:0] alpha387_2_x_locator2;
  wire [9:0] alpha387_3_x_locator3;
  wire [9:0] alpha388_0_x_locator0;
  wire [9:0] alpha388_1_x_locator1;
  wire [9:0] alpha388_2_x_locator2;
  wire [9:0] alpha388_3_x_locator3;
  wire [9:0] alpha389_0_x_locator0;
  wire [9:0] alpha389_1_x_locator1;
  wire [9:0] alpha389_2_x_locator2;
  wire [9:0] alpha389_3_x_locator3;
  wire [9:0] alpha390_0_x_locator0;
  wire [9:0] alpha390_1_x_locator1;
  wire [9:0] alpha390_2_x_locator2;
  wire [9:0] alpha390_3_x_locator3;
  wire [9:0] alpha391_0_x_locator0;
  wire [9:0] alpha391_1_x_locator1;
  wire [9:0] alpha391_2_x_locator2;
  wire [9:0] alpha391_3_x_locator3;
  wire [9:0] alpha392_0_x_locator0;
  wire [9:0] alpha392_1_x_locator1;
  wire [9:0] alpha392_2_x_locator2;
  wire [9:0] alpha392_3_x_locator3;
  wire [9:0] alpha393_0_x_locator0;
  wire [9:0] alpha393_1_x_locator1;
  wire [9:0] alpha393_2_x_locator2;
  wire [9:0] alpha393_3_x_locator3;
  wire [9:0] alpha394_0_x_locator0;
  wire [9:0] alpha394_1_x_locator1;
  wire [9:0] alpha394_2_x_locator2;
  wire [9:0] alpha394_3_x_locator3;
  wire [9:0] alpha395_0_x_locator0;
  wire [9:0] alpha395_1_x_locator1;
  wire [9:0] alpha395_2_x_locator2;
  wire [9:0] alpha395_3_x_locator3;
  wire [9:0] alpha396_0_x_locator0;
  wire [9:0] alpha396_1_x_locator1;
  wire [9:0] alpha396_2_x_locator2;
  wire [9:0] alpha396_3_x_locator3;
  wire [9:0] alpha397_0_x_locator0;
  wire [9:0] alpha397_1_x_locator1;
  wire [9:0] alpha397_2_x_locator2;
  wire [9:0] alpha397_3_x_locator3;
  wire [9:0] alpha398_0_x_locator0;
  wire [9:0] alpha398_1_x_locator1;
  wire [9:0] alpha398_2_x_locator2;
  wire [9:0] alpha398_3_x_locator3;
  wire [9:0] alpha399_0_x_locator0;
  wire [9:0] alpha399_1_x_locator1;
  wire [9:0] alpha399_2_x_locator2;
  wire [9:0] alpha399_3_x_locator3;
  wire [9:0] alpha400_0_x_locator0;
  wire [9:0] alpha400_1_x_locator1;
  wire [9:0] alpha400_2_x_locator2;
  wire [9:0] alpha400_3_x_locator3;
  wire [9:0] alpha401_0_x_locator0;
  wire [9:0] alpha401_1_x_locator1;
  wire [9:0] alpha401_2_x_locator2;
  wire [9:0] alpha401_3_x_locator3;
  wire [9:0] alpha402_0_x_locator0;
  wire [9:0] alpha402_1_x_locator1;
  wire [9:0] alpha402_2_x_locator2;
  wire [9:0] alpha402_3_x_locator3;
  wire [9:0] alpha403_0_x_locator0;
  wire [9:0] alpha403_1_x_locator1;
  wire [9:0] alpha403_2_x_locator2;
  wire [9:0] alpha403_3_x_locator3;
  wire [9:0] alpha404_0_x_locator0;
  wire [9:0] alpha404_1_x_locator1;
  wire [9:0] alpha404_2_x_locator2;
  wire [9:0] alpha404_3_x_locator3;
  wire [9:0] alpha405_0_x_locator0;
  wire [9:0] alpha405_1_x_locator1;
  wire [9:0] alpha405_2_x_locator2;
  wire [9:0] alpha405_3_x_locator3;
  wire [9:0] alpha406_0_x_locator0;
  wire [9:0] alpha406_1_x_locator1;
  wire [9:0] alpha406_2_x_locator2;
  wire [9:0] alpha406_3_x_locator3;
  wire [9:0] alpha407_0_x_locator0;
  wire [9:0] alpha407_1_x_locator1;
  wire [9:0] alpha407_2_x_locator2;
  wire [9:0] alpha407_3_x_locator3;
  wire [9:0] alpha408_0_x_locator0;
  wire [9:0] alpha408_1_x_locator1;
  wire [9:0] alpha408_2_x_locator2;
  wire [9:0] alpha408_3_x_locator3;
  wire [9:0] alpha409_0_x_locator0;
  wire [9:0] alpha409_1_x_locator1;
  wire [9:0] alpha409_2_x_locator2;
  wire [9:0] alpha409_3_x_locator3;
  wire [9:0] alpha410_0_x_locator0;
  wire [9:0] alpha410_1_x_locator1;
  wire [9:0] alpha410_2_x_locator2;
  wire [9:0] alpha410_3_x_locator3;
  wire [9:0] alpha411_0_x_locator0;
  wire [9:0] alpha411_1_x_locator1;
  wire [9:0] alpha411_2_x_locator2;
  wire [9:0] alpha411_3_x_locator3;
  wire [9:0] alpha412_0_x_locator0;
  wire [9:0] alpha412_1_x_locator1;
  wire [9:0] alpha412_2_x_locator2;
  wire [9:0] alpha412_3_x_locator3;
  wire [9:0] alpha413_0_x_locator0;
  wire [9:0] alpha413_1_x_locator1;
  wire [9:0] alpha413_2_x_locator2;
  wire [9:0] alpha413_3_x_locator3;
  wire [9:0] alpha414_0_x_locator0;
  wire [9:0] alpha414_1_x_locator1;
  wire [9:0] alpha414_2_x_locator2;
  wire [9:0] alpha414_3_x_locator3;
  wire [9:0] alpha415_0_x_locator0;
  wire [9:0] alpha415_1_x_locator1;
  wire [9:0] alpha415_2_x_locator2;
  wire [9:0] alpha415_3_x_locator3;
  wire [9:0] alpha416_0_x_locator0;
  wire [9:0] alpha416_1_x_locator1;
  wire [9:0] alpha416_2_x_locator2;
  wire [9:0] alpha416_3_x_locator3;
  wire [9:0] alpha417_0_x_locator0;
  wire [9:0] alpha417_1_x_locator1;
  wire [9:0] alpha417_2_x_locator2;
  wire [9:0] alpha417_3_x_locator3;
  wire [9:0] alpha418_0_x_locator0;
  wire [9:0] alpha418_1_x_locator1;
  wire [9:0] alpha418_2_x_locator2;
  wire [9:0] alpha418_3_x_locator3;
  wire [9:0] alpha419_0_x_locator0;
  wire [9:0] alpha419_1_x_locator1;
  wire [9:0] alpha419_2_x_locator2;
  wire [9:0] alpha419_3_x_locator3;
  wire [9:0] alpha420_0_x_locator0;
  wire [9:0] alpha420_1_x_locator1;
  wire [9:0] alpha420_2_x_locator2;
  wire [9:0] alpha420_3_x_locator3;
  wire [9:0] alpha421_0_x_locator0;
  wire [9:0] alpha421_1_x_locator1;
  wire [9:0] alpha421_2_x_locator2;
  wire [9:0] alpha421_3_x_locator3;
  wire [9:0] alpha422_0_x_locator0;
  wire [9:0] alpha422_1_x_locator1;
  wire [9:0] alpha422_2_x_locator2;
  wire [9:0] alpha422_3_x_locator3;
  wire [9:0] alpha423_0_x_locator0;
  wire [9:0] alpha423_1_x_locator1;
  wire [9:0] alpha423_2_x_locator2;
  wire [9:0] alpha423_3_x_locator3;
  wire [9:0] alpha424_0_x_locator0;
  wire [9:0] alpha424_1_x_locator1;
  wire [9:0] alpha424_2_x_locator2;
  wire [9:0] alpha424_3_x_locator3;
  wire [9:0] alpha425_0_x_locator0;
  wire [9:0] alpha425_1_x_locator1;
  wire [9:0] alpha425_2_x_locator2;
  wire [9:0] alpha425_3_x_locator3;
  wire [9:0] alpha426_0_x_locator0;
  wire [9:0] alpha426_1_x_locator1;
  wire [9:0] alpha426_2_x_locator2;
  wire [9:0] alpha426_3_x_locator3;
  wire [9:0] alpha427_0_x_locator0;
  wire [9:0] alpha427_1_x_locator1;
  wire [9:0] alpha427_2_x_locator2;
  wire [9:0] alpha427_3_x_locator3;
  wire [9:0] alpha428_0_x_locator0;
  wire [9:0] alpha428_1_x_locator1;
  wire [9:0] alpha428_2_x_locator2;
  wire [9:0] alpha428_3_x_locator3;
  wire [9:0] alpha429_0_x_locator0;
  wire [9:0] alpha429_1_x_locator1;
  wire [9:0] alpha429_2_x_locator2;
  wire [9:0] alpha429_3_x_locator3;
  wire [9:0] alpha430_0_x_locator0;
  wire [9:0] alpha430_1_x_locator1;
  wire [9:0] alpha430_2_x_locator2;
  wire [9:0] alpha430_3_x_locator3;
  wire [9:0] alpha431_0_x_locator0;
  wire [9:0] alpha431_1_x_locator1;
  wire [9:0] alpha431_2_x_locator2;
  wire [9:0] alpha431_3_x_locator3;
  wire [9:0] alpha432_0_x_locator0;
  wire [9:0] alpha432_1_x_locator1;
  wire [9:0] alpha432_2_x_locator2;
  wire [9:0] alpha432_3_x_locator3;
  wire [9:0] alpha433_0_x_locator0;
  wire [9:0] alpha433_1_x_locator1;
  wire [9:0] alpha433_2_x_locator2;
  wire [9:0] alpha433_3_x_locator3;
  wire [9:0] alpha434_0_x_locator0;
  wire [9:0] alpha434_1_x_locator1;
  wire [9:0] alpha434_2_x_locator2;
  wire [9:0] alpha434_3_x_locator3;
  wire [9:0] alpha435_0_x_locator0;
  wire [9:0] alpha435_1_x_locator1;
  wire [9:0] alpha435_2_x_locator2;
  wire [9:0] alpha435_3_x_locator3;
  wire [9:0] alpha436_0_x_locator0;
  wire [9:0] alpha436_1_x_locator1;
  wire [9:0] alpha436_2_x_locator2;
  wire [9:0] alpha436_3_x_locator3;
  wire [9:0] alpha437_0_x_locator0;
  wire [9:0] alpha437_1_x_locator1;
  wire [9:0] alpha437_2_x_locator2;
  wire [9:0] alpha437_3_x_locator3;
  wire [9:0] alpha438_0_x_locator0;
  wire [9:0] alpha438_1_x_locator1;
  wire [9:0] alpha438_2_x_locator2;
  wire [9:0] alpha438_3_x_locator3;
  wire [9:0] alpha439_0_x_locator0;
  wire [9:0] alpha439_1_x_locator1;
  wire [9:0] alpha439_2_x_locator2;
  wire [9:0] alpha439_3_x_locator3;
  wire [9:0] alpha440_0_x_locator0;
  wire [9:0] alpha440_1_x_locator1;
  wire [9:0] alpha440_2_x_locator2;
  wire [9:0] alpha440_3_x_locator3;
  wire [9:0] alpha441_0_x_locator0;
  wire [9:0] alpha441_1_x_locator1;
  wire [9:0] alpha441_2_x_locator2;
  wire [9:0] alpha441_3_x_locator3;
  wire [9:0] alpha442_0_x_locator0;
  wire [9:0] alpha442_1_x_locator1;
  wire [9:0] alpha442_2_x_locator2;
  wire [9:0] alpha442_3_x_locator3;
  wire [9:0] alpha443_0_x_locator0;
  wire [9:0] alpha443_1_x_locator1;
  wire [9:0] alpha443_2_x_locator2;
  wire [9:0] alpha443_3_x_locator3;
  wire [9:0] alpha444_0_x_locator0;
  wire [9:0] alpha444_1_x_locator1;
  wire [9:0] alpha444_2_x_locator2;
  wire [9:0] alpha444_3_x_locator3;
  wire [9:0] alpha445_0_x_locator0;
  wire [9:0] alpha445_1_x_locator1;
  wire [9:0] alpha445_2_x_locator2;
  wire [9:0] alpha445_3_x_locator3;
  wire [9:0] alpha446_0_x_locator0;
  wire [9:0] alpha446_1_x_locator1;
  wire [9:0] alpha446_2_x_locator2;
  wire [9:0] alpha446_3_x_locator3;
  wire [9:0] alpha447_0_x_locator0;
  wire [9:0] alpha447_1_x_locator1;
  wire [9:0] alpha447_2_x_locator2;
  wire [9:0] alpha447_3_x_locator3;
  wire [9:0] alpha448_0_x_locator0;
  wire [9:0] alpha448_1_x_locator1;
  wire [9:0] alpha448_2_x_locator2;
  wire [9:0] alpha448_3_x_locator3;
  wire [9:0] alpha449_0_x_locator0;
  wire [9:0] alpha449_1_x_locator1;
  wire [9:0] alpha449_2_x_locator2;
  wire [9:0] alpha449_3_x_locator3;
  wire [9:0] alpha450_0_x_locator0;
  wire [9:0] alpha450_1_x_locator1;
  wire [9:0] alpha450_2_x_locator2;
  wire [9:0] alpha450_3_x_locator3;
  wire [9:0] alpha451_0_x_locator0;
  wire [9:0] alpha451_1_x_locator1;
  wire [9:0] alpha451_2_x_locator2;
  wire [9:0] alpha451_3_x_locator3;
  wire [9:0] alpha452_0_x_locator0;
  wire [9:0] alpha452_1_x_locator1;
  wire [9:0] alpha452_2_x_locator2;
  wire [9:0] alpha452_3_x_locator3;
  wire [9:0] alpha453_0_x_locator0;
  wire [9:0] alpha453_1_x_locator1;
  wire [9:0] alpha453_2_x_locator2;
  wire [9:0] alpha453_3_x_locator3;
  wire [9:0] alpha454_0_x_locator0;
  wire [9:0] alpha454_1_x_locator1;
  wire [9:0] alpha454_2_x_locator2;
  wire [9:0] alpha454_3_x_locator3;
  wire [9:0] alpha455_0_x_locator0;
  wire [9:0] alpha455_1_x_locator1;
  wire [9:0] alpha455_2_x_locator2;
  wire [9:0] alpha455_3_x_locator3;
  wire [9:0] alpha456_0_x_locator0;
  wire [9:0] alpha456_1_x_locator1;
  wire [9:0] alpha456_2_x_locator2;
  wire [9:0] alpha456_3_x_locator3;
  wire [9:0] alpha457_0_x_locator0;
  wire [9:0] alpha457_1_x_locator1;
  wire [9:0] alpha457_2_x_locator2;
  wire [9:0] alpha457_3_x_locator3;
  wire [9:0] alpha458_0_x_locator0;
  wire [9:0] alpha458_1_x_locator1;
  wire [9:0] alpha458_2_x_locator2;
  wire [9:0] alpha458_3_x_locator3;
  wire [9:0] alpha459_0_x_locator0;
  wire [9:0] alpha459_1_x_locator1;
  wire [9:0] alpha459_2_x_locator2;
  wire [9:0] alpha459_3_x_locator3;
  wire [9:0] alpha460_0_x_locator0;
  wire [9:0] alpha460_1_x_locator1;
  wire [9:0] alpha460_2_x_locator2;
  wire [9:0] alpha460_3_x_locator3;
  wire [9:0] alpha461_0_x_locator0;
  wire [9:0] alpha461_1_x_locator1;
  wire [9:0] alpha461_2_x_locator2;
  wire [9:0] alpha461_3_x_locator3;
  wire [9:0] alpha462_0_x_locator0;
  wire [9:0] alpha462_1_x_locator1;
  wire [9:0] alpha462_2_x_locator2;
  wire [9:0] alpha462_3_x_locator3;
  wire [9:0] alpha463_0_x_locator0;
  wire [9:0] alpha463_1_x_locator1;
  wire [9:0] alpha463_2_x_locator2;
  wire [9:0] alpha463_3_x_locator3;
  wire [9:0] alpha464_0_x_locator0;
  wire [9:0] alpha464_1_x_locator1;
  wire [9:0] alpha464_2_x_locator2;
  wire [9:0] alpha464_3_x_locator3;
  wire [9:0] alpha465_0_x_locator0;
  wire [9:0] alpha465_1_x_locator1;
  wire [9:0] alpha465_2_x_locator2;
  wire [9:0] alpha465_3_x_locator3;
  wire [9:0] alpha466_0_x_locator0;
  wire [9:0] alpha466_1_x_locator1;
  wire [9:0] alpha466_2_x_locator2;
  wire [9:0] alpha466_3_x_locator3;
  wire [9:0] alpha467_0_x_locator0;
  wire [9:0] alpha467_1_x_locator1;
  wire [9:0] alpha467_2_x_locator2;
  wire [9:0] alpha467_3_x_locator3;
  wire [9:0] alpha468_0_x_locator0;
  wire [9:0] alpha468_1_x_locator1;
  wire [9:0] alpha468_2_x_locator2;
  wire [9:0] alpha468_3_x_locator3;
  wire [9:0] alpha469_0_x_locator0;
  wire [9:0] alpha469_1_x_locator1;
  wire [9:0] alpha469_2_x_locator2;
  wire [9:0] alpha469_3_x_locator3;
  wire [9:0] alpha470_0_x_locator0;
  wire [9:0] alpha470_1_x_locator1;
  wire [9:0] alpha470_2_x_locator2;
  wire [9:0] alpha470_3_x_locator3;
  wire [9:0] alpha471_0_x_locator0;
  wire [9:0] alpha471_1_x_locator1;
  wire [9:0] alpha471_2_x_locator2;
  wire [9:0] alpha471_3_x_locator3;
  wire [9:0] alpha472_0_x_locator0;
  wire [9:0] alpha472_1_x_locator1;
  wire [9:0] alpha472_2_x_locator2;
  wire [9:0] alpha472_3_x_locator3;
  wire [9:0] alpha473_0_x_locator0;
  wire [9:0] alpha473_1_x_locator1;
  wire [9:0] alpha473_2_x_locator2;
  wire [9:0] alpha473_3_x_locator3;
  wire [9:0] alpha474_0_x_locator0;
  wire [9:0] alpha474_1_x_locator1;
  wire [9:0] alpha474_2_x_locator2;
  wire [9:0] alpha474_3_x_locator3;
  wire [9:0] alpha475_0_x_locator0;
  wire [9:0] alpha475_1_x_locator1;
  wire [9:0] alpha475_2_x_locator2;
  wire [9:0] alpha475_3_x_locator3;
  wire [9:0] alpha476_0_x_locator0;
  wire [9:0] alpha476_1_x_locator1;
  wire [9:0] alpha476_2_x_locator2;
  wire [9:0] alpha476_3_x_locator3;
  wire [9:0] alpha477_0_x_locator0;
  wire [9:0] alpha477_1_x_locator1;
  wire [9:0] alpha477_2_x_locator2;
  wire [9:0] alpha477_3_x_locator3;
  wire [9:0] alpha478_0_x_locator0;
  wire [9:0] alpha478_1_x_locator1;
  wire [9:0] alpha478_2_x_locator2;
  wire [9:0] alpha478_3_x_locator3;
  wire [9:0] alpha479_0_x_locator0;
  wire [9:0] alpha479_1_x_locator1;
  wire [9:0] alpha479_2_x_locator2;
  wire [9:0] alpha479_3_x_locator3;
  wire [9:0] alpha480_0_x_locator0;
  wire [9:0] alpha480_1_x_locator1;
  wire [9:0] alpha480_2_x_locator2;
  wire [9:0] alpha480_3_x_locator3;
  wire [9:0] alpha481_0_x_locator0;
  wire [9:0] alpha481_1_x_locator1;
  wire [9:0] alpha481_2_x_locator2;
  wire [9:0] alpha481_3_x_locator3;
  wire [9:0] alpha482_0_x_locator0;
  wire [9:0] alpha482_1_x_locator1;
  wire [9:0] alpha482_2_x_locator2;
  wire [9:0] alpha482_3_x_locator3;
  wire [9:0] alpha483_0_x_locator0;
  wire [9:0] alpha483_1_x_locator1;
  wire [9:0] alpha483_2_x_locator2;
  wire [9:0] alpha483_3_x_locator3;
  wire [9:0] alpha484_0_x_locator0;
  wire [9:0] alpha484_1_x_locator1;
  wire [9:0] alpha484_2_x_locator2;
  wire [9:0] alpha484_3_x_locator3;
  wire [9:0] alpha485_0_x_locator0;
  wire [9:0] alpha485_1_x_locator1;
  wire [9:0] alpha485_2_x_locator2;
  wire [9:0] alpha485_3_x_locator3;
  wire [9:0] alpha486_0_x_locator0;
  wire [9:0] alpha486_1_x_locator1;
  wire [9:0] alpha486_2_x_locator2;
  wire [9:0] alpha486_3_x_locator3;
  wire [9:0] alpha487_0_x_locator0;
  wire [9:0] alpha487_1_x_locator1;
  wire [9:0] alpha487_2_x_locator2;
  wire [9:0] alpha487_3_x_locator3;
  wire [9:0] alpha488_0_x_locator0;
  wire [9:0] alpha488_1_x_locator1;
  wire [9:0] alpha488_2_x_locator2;
  wire [9:0] alpha488_3_x_locator3;
  wire [9:0] alpha489_0_x_locator0;
  wire [9:0] alpha489_1_x_locator1;
  wire [9:0] alpha489_2_x_locator2;
  wire [9:0] alpha489_3_x_locator3;
  wire [9:0] alpha490_0_x_locator0;
  wire [9:0] alpha490_1_x_locator1;
  wire [9:0] alpha490_2_x_locator2;
  wire [9:0] alpha490_3_x_locator3;
  wire [9:0] alpha491_0_x_locator0;
  wire [9:0] alpha491_1_x_locator1;
  wire [9:0] alpha491_2_x_locator2;
  wire [9:0] alpha491_3_x_locator3;
  wire [9:0] alpha492_0_x_locator0;
  wire [9:0] alpha492_1_x_locator1;
  wire [9:0] alpha492_2_x_locator2;
  wire [9:0] alpha492_3_x_locator3;
  wire [9:0] alpha493_0_x_locator0;
  wire [9:0] alpha493_1_x_locator1;
  wire [9:0] alpha493_2_x_locator2;
  wire [9:0] alpha493_3_x_locator3;
  wire [9:0] alpha494_0_x_locator0;
  wire [9:0] alpha494_1_x_locator1;
  wire [9:0] alpha494_2_x_locator2;
  wire [9:0] alpha494_3_x_locator3;
  wire [9:0] alpha495_0_x_locator0;
  wire [9:0] alpha495_1_x_locator1;
  wire [9:0] alpha495_2_x_locator2;
  wire [9:0] alpha495_3_x_locator3;
  wire [9:0] alpha496_0_x_locator0;
  wire [9:0] alpha496_1_x_locator1;
  wire [9:0] alpha496_2_x_locator2;
  wire [9:0] alpha496_3_x_locator3;
  wire [9:0] alpha497_0_x_locator0;
  wire [9:0] alpha497_1_x_locator1;
  wire [9:0] alpha497_2_x_locator2;
  wire [9:0] alpha497_3_x_locator3;
  wire [9:0] alpha498_0_x_locator0;
  wire [9:0] alpha498_1_x_locator1;
  wire [9:0] alpha498_2_x_locator2;
  wire [9:0] alpha498_3_x_locator3;
  wire [9:0] alpha499_0_x_locator0;
  wire [9:0] alpha499_1_x_locator1;
  wire [9:0] alpha499_2_x_locator2;
  wire [9:0] alpha499_3_x_locator3;
  wire [9:0] alpha500_0_x_locator0;
  wire [9:0] alpha500_1_x_locator1;
  wire [9:0] alpha500_2_x_locator2;
  wire [9:0] alpha500_3_x_locator3;
  wire [9:0] alpha501_0_x_locator0;
  wire [9:0] alpha501_1_x_locator1;
  wire [9:0] alpha501_2_x_locator2;
  wire [9:0] alpha501_3_x_locator3;
  wire [9:0] alpha502_0_x_locator0;
  wire [9:0] alpha502_1_x_locator1;
  wire [9:0] alpha502_2_x_locator2;
  wire [9:0] alpha502_3_x_locator3;
  wire [9:0] alpha503_0_x_locator0;
  wire [9:0] alpha503_1_x_locator1;
  wire [9:0] alpha503_2_x_locator2;
  wire [9:0] alpha503_3_x_locator3;
  wire [9:0] alpha504_0_x_locator0;
  wire [9:0] alpha504_1_x_locator1;
  wire [9:0] alpha504_2_x_locator2;
  wire [9:0] alpha504_3_x_locator3;
  wire [9:0] alpha505_0_x_locator0;
  wire [9:0] alpha505_1_x_locator1;
  wire [9:0] alpha505_2_x_locator2;
  wire [9:0] alpha505_3_x_locator3;
  wire [9:0] alpha506_0_x_locator0;
  wire [9:0] alpha506_1_x_locator1;
  wire [9:0] alpha506_2_x_locator2;
  wire [9:0] alpha506_3_x_locator3;
  wire [9:0] alpha507_0_x_locator0;
  wire [9:0] alpha507_1_x_locator1;
  wire [9:0] alpha507_2_x_locator2;
  wire [9:0] alpha507_3_x_locator3;
  wire [9:0] alpha508_0_x_locator0;
  wire [9:0] alpha508_1_x_locator1;
  wire [9:0] alpha508_2_x_locator2;
  wire [9:0] alpha508_3_x_locator3;
  wire [9:0] alpha509_0_x_locator0;
  wire [9:0] alpha509_1_x_locator1;
  wire [9:0] alpha509_2_x_locator2;
  wire [9:0] alpha509_3_x_locator3;
  wire [9:0] alpha510_0_x_locator0;
  wire [9:0] alpha510_1_x_locator1;
  wire [9:0] alpha510_2_x_locator2;
  wire [9:0] alpha510_3_x_locator3;
  wire [9:0] alpha511_0_x_locator0;
  wire [9:0] alpha511_1_x_locator1;
  wire [9:0] alpha511_2_x_locator2;
  wire [9:0] alpha511_3_x_locator3;
  wire [9:0] alpha512_0_x_locator0;
  wire [9:0] alpha512_1_x_locator1;
  wire [9:0] alpha512_2_x_locator2;
  wire [9:0] alpha512_3_x_locator3;
  wire [9:0] alpha513_0_x_locator0;
  wire [9:0] alpha513_1_x_locator1;
  wire [9:0] alpha513_2_x_locator2;
  wire [9:0] alpha513_3_x_locator3;
  wire [9:0] alpha514_0_x_locator0;
  wire [9:0] alpha514_1_x_locator1;
  wire [9:0] alpha514_2_x_locator2;
  wire [9:0] alpha514_3_x_locator3;
  wire [9:0] alpha515_0_x_locator0;
  wire [9:0] alpha515_1_x_locator1;
  wire [9:0] alpha515_2_x_locator2;
  wire [9:0] alpha515_3_x_locator3;
  wire [9:0] alpha516_0_x_locator0;
  wire [9:0] alpha516_1_x_locator1;
  wire [9:0] alpha516_2_x_locator2;
  wire [9:0] alpha516_3_x_locator3;
  wire [9:0] alpha517_0_x_locator0;
  wire [9:0] alpha517_1_x_locator1;
  wire [9:0] alpha517_2_x_locator2;
  wire [9:0] alpha517_3_x_locator3;
  wire [9:0] alpha518_0_x_locator0;
  wire [9:0] alpha518_1_x_locator1;
  wire [9:0] alpha518_2_x_locator2;
  wire [9:0] alpha518_3_x_locator3;
  wire [9:0] alpha519_0_x_locator0;
  wire [9:0] alpha519_1_x_locator1;
  wire [9:0] alpha519_2_x_locator2;
  wire [9:0] alpha519_3_x_locator3;
  wire [9:0] alpha520_0_x_locator0;
  wire [9:0] alpha520_1_x_locator1;
  wire [9:0] alpha520_2_x_locator2;
  wire [9:0] alpha520_3_x_locator3;
  wire [9:0] alpha521_0_x_locator0;
  wire [9:0] alpha521_1_x_locator1;
  wire [9:0] alpha521_2_x_locator2;
  wire [9:0] alpha521_3_x_locator3;
  wire [9:0] alpha522_0_x_locator0;
  wire [9:0] alpha522_1_x_locator1;
  wire [9:0] alpha522_2_x_locator2;
  wire [9:0] alpha522_3_x_locator3;
  wire [9:0] alpha523_0_x_locator0;
  wire [9:0] alpha523_1_x_locator1;
  wire [9:0] alpha523_2_x_locator2;
  wire [9:0] alpha523_3_x_locator3;
  wire [9:0] alpha524_0_x_locator0;
  wire [9:0] alpha524_1_x_locator1;
  wire [9:0] alpha524_2_x_locator2;
  wire [9:0] alpha524_3_x_locator3;
  wire [9:0] alpha525_0_x_locator0;
  wire [9:0] alpha525_1_x_locator1;
  wire [9:0] alpha525_2_x_locator2;
  wire [9:0] alpha525_3_x_locator3;
  wire [9:0] alpha526_0_x_locator0;
  wire [9:0] alpha526_1_x_locator1;
  wire [9:0] alpha526_2_x_locator2;
  wire [9:0] alpha526_3_x_locator3;
  wire [9:0] alpha527_0_x_locator0;
  wire [9:0] alpha527_1_x_locator1;
  wire [9:0] alpha527_2_x_locator2;
  wire [9:0] alpha527_3_x_locator3;
  wire [9:0] alpha528_0_x_locator0;
  wire [9:0] alpha528_1_x_locator1;
  wire [9:0] alpha528_2_x_locator2;
  wire [9:0] alpha528_3_x_locator3;
  wire [9:0] alpha529_0_x_locator0;
  wire [9:0] alpha529_1_x_locator1;
  wire [9:0] alpha529_2_x_locator2;
  wire [9:0] alpha529_3_x_locator3;
  wire [9:0] alpha530_0_x_locator0;
  wire [9:0] alpha530_1_x_locator1;
  wire [9:0] alpha530_2_x_locator2;
  wire [9:0] alpha530_3_x_locator3;
  wire [9:0] alpha531_0_x_locator0;
  wire [9:0] alpha531_1_x_locator1;
  wire [9:0] alpha531_2_x_locator2;
  wire [9:0] alpha531_3_x_locator3;
  wire [9:0] alpha532_0_x_locator0;
  wire [9:0] alpha532_1_x_locator1;
  wire [9:0] alpha532_2_x_locator2;
  wire [9:0] alpha532_3_x_locator3;
  wire [9:0] alpha533_0_x_locator0;
  wire [9:0] alpha533_1_x_locator1;
  wire [9:0] alpha533_2_x_locator2;
  wire [9:0] alpha533_3_x_locator3;
  wire [9:0] alpha534_0_x_locator0;
  wire [9:0] alpha534_1_x_locator1;
  wire [9:0] alpha534_2_x_locator2;
  wire [9:0] alpha534_3_x_locator3;
  wire [9:0] alpha535_0_x_locator0;
  wire [9:0] alpha535_1_x_locator1;
  wire [9:0] alpha535_2_x_locator2;
  wire [9:0] alpha535_3_x_locator3;
  wire [9:0] alpha536_0_x_locator0;
  wire [9:0] alpha536_1_x_locator1;
  wire [9:0] alpha536_2_x_locator2;
  wire [9:0] alpha536_3_x_locator3;
  wire [9:0] alpha537_0_x_locator0;
  wire [9:0] alpha537_1_x_locator1;
  wire [9:0] alpha537_2_x_locator2;
  wire [9:0] alpha537_3_x_locator3;
  wire [9:0] alpha538_0_x_locator0;
  wire [9:0] alpha538_1_x_locator1;
  wire [9:0] alpha538_2_x_locator2;
  wire [9:0] alpha538_3_x_locator3;
  wire [9:0] alpha539_0_x_locator0;
  wire [9:0] alpha539_1_x_locator1;
  wire [9:0] alpha539_2_x_locator2;
  wire [9:0] alpha539_3_x_locator3;
  wire [9:0] alpha540_0_x_locator0;
  wire [9:0] alpha540_1_x_locator1;
  wire [9:0] alpha540_2_x_locator2;
  wire [9:0] alpha540_3_x_locator3;
  wire [9:0] alpha541_0_x_locator0;
  wire [9:0] alpha541_1_x_locator1;
  wire [9:0] alpha541_2_x_locator2;
  wire [9:0] alpha541_3_x_locator3;

  gfmult gfm_alpha0_0_x_locator0(10'b0000000001, locator0, alpha0_0_x_locator0);
  gfmult gfm_alpha0_1_x_locator1(10'b0000000001, locator1, alpha0_1_x_locator1);
  gfmult gfm_alpha0_2_x_locator2(10'b0000000001, locator2, alpha0_2_x_locator2);
  gfmult gfm_alpha0_3_x_locator3(10'b0000000001, locator3, alpha0_3_x_locator3);
  gfmult gfm_alpha1_0_x_locator0(10'b0000000001, locator0, alpha1_0_x_locator0);
  gfmult gfm_alpha1_1_x_locator1(10'b1000000100, locator1, alpha1_1_x_locator1);
  gfmult gfm_alpha1_2_x_locator2(10'b0100000010, locator2, alpha1_2_x_locator2);
  gfmult gfm_alpha1_3_x_locator3(10'b0010000001, locator3, alpha1_3_x_locator3);
  gfmult gfm_alpha2_0_x_locator0(10'b0000000001, locator0, alpha2_0_x_locator0);
  gfmult gfm_alpha2_1_x_locator1(10'b0100000010, locator1, alpha2_1_x_locator1);
  gfmult gfm_alpha2_2_x_locator2(10'b1001000100, locator2, alpha2_2_x_locator2);
  gfmult gfm_alpha2_3_x_locator3(10'b0010010001, locator3, alpha2_3_x_locator3);
  gfmult gfm_alpha3_0_x_locator0(10'b0000000001, locator0, alpha3_0_x_locator0);
  gfmult gfm_alpha3_1_x_locator1(10'b0010000001, locator1, alpha3_1_x_locator1);
  gfmult gfm_alpha3_2_x_locator2(10'b0010010001, locator2, alpha3_2_x_locator2);
  gfmult gfm_alpha3_3_x_locator3(10'b0010010011, locator3, alpha3_3_x_locator3);
  gfmult gfm_alpha4_0_x_locator0(10'b0000000001, locator0, alpha4_0_x_locator0);
  gfmult gfm_alpha4_1_x_locator1(10'b1001000100, locator1, alpha4_1_x_locator1);
  gfmult gfm_alpha4_2_x_locator2(10'b0100100110, locator2, alpha4_2_x_locator2);
  gfmult gfm_alpha4_3_x_locator3(10'b0110010001, locator3, alpha4_3_x_locator3);
  gfmult gfm_alpha5_0_x_locator0(10'b0000000001, locator0, alpha5_0_x_locator0);
  gfmult gfm_alpha5_1_x_locator1(10'b0100100010, locator1, alpha5_1_x_locator1);
  gfmult gfm_alpha5_2_x_locator2(10'b1001001101, locator2, alpha5_2_x_locator2);
  gfmult gfm_alpha5_3_x_locator3(10'b0010110011, locator3, alpha5_3_x_locator3);
  gfmult gfm_alpha6_0_x_locator0(10'b0000000001, locator0, alpha6_0_x_locator0);
  gfmult gfm_alpha6_1_x_locator1(10'b0010010001, locator1, alpha6_1_x_locator1);
  gfmult gfm_alpha6_2_x_locator2(10'b0110010001, locator2, alpha6_2_x_locator2);
  gfmult gfm_alpha6_3_x_locator3(10'b0110010101, locator3, alpha6_3_x_locator3);
  gfmult gfm_alpha7_0_x_locator0(10'b0000000001, locator0, alpha7_0_x_locator0);
  gfmult gfm_alpha7_1_x_locator1(10'b1001001100, locator1, alpha7_1_x_locator1);
  gfmult gfm_alpha7_2_x_locator2(10'b0101100110, locator2, alpha7_2_x_locator2);
  gfmult gfm_alpha7_3_x_locator3(10'b1010110111, locator3, alpha7_3_x_locator3);
  gfmult gfm_alpha8_0_x_locator0(10'b0000000001, locator0, alpha8_0_x_locator0);
  gfmult gfm_alpha8_1_x_locator1(10'b0100100110, locator1, alpha8_1_x_locator1);
  gfmult gfm_alpha8_2_x_locator2(10'b1001011101, locator2, alpha8_2_x_locator2);
  gfmult gfm_alpha8_3_x_locator3(10'b1111010001, locator3, alpha8_3_x_locator3);
  gfmult gfm_alpha9_0_x_locator0(10'b0000000001, locator0, alpha9_0_x_locator0);
  gfmult gfm_alpha9_1_x_locator1(10'b0010010011, locator1, alpha9_1_x_locator1);
  gfmult gfm_alpha9_2_x_locator2(10'b0110010101, locator2, alpha9_2_x_locator2);
  gfmult gfm_alpha9_3_x_locator3(10'b0011111011, locator3, alpha9_3_x_locator3);
  gfmult gfm_alpha10_0_x_locator0(10'b0000000001, locator0, alpha10_0_x_locator0);
  gfmult gfm_alpha10_1_x_locator1(10'b1001001101, locator1, alpha10_1_x_locator1);
  gfmult gfm_alpha10_2_x_locator2(10'b0101100111, locator2, alpha10_2_x_locator2);
  gfmult gfm_alpha10_3_x_locator3(10'b0110011100, locator3, alpha10_3_x_locator3);
  gfmult gfm_alpha11_0_x_locator0(10'b0000000001, locator0, alpha11_0_x_locator0);
  gfmult gfm_alpha11_1_x_locator1(10'b1100100010, locator1, alpha11_1_x_locator1);
  gfmult gfm_alpha11_2_x_locator2(10'b1101011111, locator2, alpha11_2_x_locator2);
  gfmult gfm_alpha11_3_x_locator3(10'b1000110111, locator3, alpha11_3_x_locator3);
  gfmult gfm_alpha12_0_x_locator0(10'b0000000001, locator0, alpha12_0_x_locator0);
  gfmult gfm_alpha12_1_x_locator1(10'b0110010001, locator1, alpha12_1_x_locator1);
  gfmult gfm_alpha12_2_x_locator2(10'b1111010001, locator2, alpha12_2_x_locator2);
  gfmult gfm_alpha12_3_x_locator3(10'b1111000001, locator3, alpha12_3_x_locator3);
  gfmult gfm_alpha13_0_x_locator0(10'b0000000001, locator0, alpha13_0_x_locator0);
  gfmult gfm_alpha13_1_x_locator1(10'b1011001100, locator1, alpha13_1_x_locator1);
  gfmult gfm_alpha13_2_x_locator2(10'b0111110110, locator2, alpha13_2_x_locator2);
  gfmult gfm_alpha13_3_x_locator3(10'b0011111001, locator3, alpha13_3_x_locator3);
  gfmult gfm_alpha14_0_x_locator0(10'b0000000001, locator0, alpha14_0_x_locator0);
  gfmult gfm_alpha14_1_x_locator1(10'b0101100110, locator1, alpha14_1_x_locator1);
  gfmult gfm_alpha14_2_x_locator2(10'b1001111001, locator2, alpha14_2_x_locator2);
  gfmult gfm_alpha14_3_x_locator3(10'b0010011110, locator3, alpha14_3_x_locator3);
  gfmult gfm_alpha15_0_x_locator0(10'b0000000001, locator0, alpha15_0_x_locator0);
  gfmult gfm_alpha15_1_x_locator1(10'b0010110011, locator1, alpha15_1_x_locator1);
  gfmult gfm_alpha15_2_x_locator2(10'b0110011100, locator2, alpha15_2_x_locator2);
  gfmult gfm_alpha15_3_x_locator3(10'b1100010101, locator3, alpha15_3_x_locator3);
  gfmult gfm_alpha16_0_x_locator0(10'b0000000001, locator0, alpha16_0_x_locator0);
  gfmult gfm_alpha16_1_x_locator1(10'b1001011101, locator1, alpha16_1_x_locator1);
  gfmult gfm_alpha16_2_x_locator2(10'b0001100111, locator2, alpha16_2_x_locator2);
  gfmult gfm_alpha16_3_x_locator3(10'b1011100111, locator3, alpha16_3_x_locator3);
  gfmult gfm_alpha17_0_x_locator0(10'b0000000001, locator0, alpha17_0_x_locator0);
  gfmult gfm_alpha17_1_x_locator1(10'b1100101010, locator1, alpha17_1_x_locator1);
  gfmult gfm_alpha17_2_x_locator2(10'b1100011111, locator2, alpha17_2_x_locator2);
  gfmult gfm_alpha17_3_x_locator3(10'b1111011011, locator3, alpha17_3_x_locator3);
  gfmult gfm_alpha18_0_x_locator0(10'b0000000001, locator0, alpha18_0_x_locator0);
  gfmult gfm_alpha18_1_x_locator1(10'b0110010101, locator1, alpha18_1_x_locator1);
  gfmult gfm_alpha18_2_x_locator2(10'b1111000001, locator2, alpha18_2_x_locator2);
  gfmult gfm_alpha18_3_x_locator3(10'b0111111000, locator3, alpha18_3_x_locator3);
  gfmult gfm_alpha19_0_x_locator0(10'b0000000001, locator0, alpha19_0_x_locator0);
  gfmult gfm_alpha19_1_x_locator1(10'b1011001110, locator1, alpha19_1_x_locator1);
  gfmult gfm_alpha19_2_x_locator2(10'b0111110010, locator2, alpha19_2_x_locator2);
  gfmult gfm_alpha19_3_x_locator3(10'b0000111111, locator3, alpha19_3_x_locator3);
  gfmult gfm_alpha20_0_x_locator0(10'b0000000001, locator0, alpha20_0_x_locator0);
  gfmult gfm_alpha20_1_x_locator1(10'b0101100111, locator1, alpha20_1_x_locator1);
  gfmult gfm_alpha20_2_x_locator2(10'b1001111000, locator2, alpha20_2_x_locator2);
  gfmult gfm_alpha20_3_x_locator3(10'b1110000000, locator3, alpha20_3_x_locator3);
  gfmult gfm_alpha21_0_x_locator0(10'b0000000001, locator0, alpha21_0_x_locator0);
  gfmult gfm_alpha21_1_x_locator1(10'b1010110111, locator1, alpha21_1_x_locator1);
  gfmult gfm_alpha21_2_x_locator2(10'b0010011110, locator2, alpha21_2_x_locator2);
  gfmult gfm_alpha21_3_x_locator3(10'b0001110000, locator3, alpha21_3_x_locator3);
  gfmult gfm_alpha22_0_x_locator0(10'b0000000001, locator0, alpha22_0_x_locator0);
  gfmult gfm_alpha22_1_x_locator1(10'b1101011111, locator1, alpha22_1_x_locator1);
  gfmult gfm_alpha22_2_x_locator2(10'b1000100011, locator2, alpha22_2_x_locator2);
  gfmult gfm_alpha22_3_x_locator3(10'b0000001110, locator3, alpha22_3_x_locator3);
  gfmult gfm_alpha23_0_x_locator0(10'b0000000001, locator0, alpha23_0_x_locator0);
  gfmult gfm_alpha23_1_x_locator1(10'b1110101011, locator1, alpha23_1_x_locator1);
  gfmult gfm_alpha23_2_x_locator2(10'b1110001110, locator2, alpha23_2_x_locator2);
  gfmult gfm_alpha23_3_x_locator3(10'b1100000111, locator3, alpha23_3_x_locator3);
  gfmult gfm_alpha24_0_x_locator0(10'b0000000001, locator0, alpha24_0_x_locator0);
  gfmult gfm_alpha24_1_x_locator1(10'b1111010001, locator1, alpha24_1_x_locator1);
  gfmult gfm_alpha24_2_x_locator2(10'b1011100111, locator2, alpha24_2_x_locator2);
  gfmult gfm_alpha24_3_x_locator3(10'b1111100111, locator3, alpha24_3_x_locator3);
  gfmult gfm_alpha25_0_x_locator0(10'b0000000001, locator0, alpha25_0_x_locator0);
  gfmult gfm_alpha25_1_x_locator1(10'b1111101100, locator1, alpha25_1_x_locator1);
  gfmult gfm_alpha25_2_x_locator2(10'b1110111111, locator2, alpha25_2_x_locator2);
  gfmult gfm_alpha25_3_x_locator3(10'b1111111011, locator3, alpha25_3_x_locator3);
  gfmult gfm_alpha26_0_x_locator0(10'b0000000001, locator0, alpha26_0_x_locator0);
  gfmult gfm_alpha26_1_x_locator1(10'b0111110110, locator1, alpha26_1_x_locator1);
  gfmult gfm_alpha26_2_x_locator2(10'b1111101001, locator2, alpha26_2_x_locator2);
  gfmult gfm_alpha26_3_x_locator3(10'b0111111100, locator3, alpha26_3_x_locator3);
  gfmult gfm_alpha27_0_x_locator0(10'b0000000001, locator0, alpha27_0_x_locator0);
  gfmult gfm_alpha27_1_x_locator1(10'b0011111011, locator1, alpha27_1_x_locator1);
  gfmult gfm_alpha27_2_x_locator2(10'b0111111000, locator2, alpha27_2_x_locator2);
  gfmult gfm_alpha27_3_x_locator3(10'b1000111011, locator3, alpha27_3_x_locator3);
  gfmult gfm_alpha28_0_x_locator0(10'b0000000001, locator0, alpha28_0_x_locator0);
  gfmult gfm_alpha28_1_x_locator1(10'b1001111001, locator1, alpha28_1_x_locator1);
  gfmult gfm_alpha28_2_x_locator2(10'b0001111110, locator2, alpha28_2_x_locator2);
  gfmult gfm_alpha28_3_x_locator3(10'b0111000100, locator3, alpha28_3_x_locator3);
  gfmult gfm_alpha29_0_x_locator0(10'b0000000001, locator0, alpha29_0_x_locator0);
  gfmult gfm_alpha29_1_x_locator1(10'b1100111000, locator1, alpha29_1_x_locator1);
  gfmult gfm_alpha29_2_x_locator2(10'b1000011011, locator2, alpha29_2_x_locator2);
  gfmult gfm_alpha29_3_x_locator3(10'b1000111100, locator3, alpha29_3_x_locator3);
  gfmult gfm_alpha30_0_x_locator0(10'b0000000001, locator0, alpha30_0_x_locator0);
  gfmult gfm_alpha30_1_x_locator1(10'b0110011100, locator1, alpha30_1_x_locator1);
  gfmult gfm_alpha30_2_x_locator2(10'b1110000000, locator2, alpha30_2_x_locator2);
  gfmult gfm_alpha30_3_x_locator3(10'b1001000011, locator3, alpha30_3_x_locator3);
  gfmult gfm_alpha31_0_x_locator0(10'b0000000001, locator0, alpha31_0_x_locator0);
  gfmult gfm_alpha31_1_x_locator1(10'b0011001110, locator1, alpha31_1_x_locator1);
  gfmult gfm_alpha31_2_x_locator2(10'b0011100000, locator2, alpha31_2_x_locator2);
  gfmult gfm_alpha31_3_x_locator3(10'b0111001011, locator3, alpha31_3_x_locator3);
  gfmult gfm_alpha32_0_x_locator0(10'b0000000001, locator0, alpha32_0_x_locator0);
  gfmult gfm_alpha32_1_x_locator1(10'b0001100111, locator1, alpha32_1_x_locator1);
  gfmult gfm_alpha32_2_x_locator2(10'b0000111000, locator2, alpha32_2_x_locator2);
  gfmult gfm_alpha32_3_x_locator3(10'b0110111010, locator3, alpha32_3_x_locator3);
  gfmult gfm_alpha33_0_x_locator0(10'b0000000001, locator0, alpha33_0_x_locator0);
  gfmult gfm_alpha33_1_x_locator1(10'b1000110111, locator1, alpha33_1_x_locator1);
  gfmult gfm_alpha33_2_x_locator2(10'b0000001110, locator2, alpha33_2_x_locator2);
  gfmult gfm_alpha33_3_x_locator3(10'b0100110101, locator3, alpha33_3_x_locator3);
  gfmult gfm_alpha34_0_x_locator0(10'b0000000001, locator0, alpha34_0_x_locator0);
  gfmult gfm_alpha34_1_x_locator1(10'b1100011111, locator1, alpha34_1_x_locator1);
  gfmult gfm_alpha34_2_x_locator2(10'b1000000111, locator2, alpha34_2_x_locator2);
  gfmult gfm_alpha34_3_x_locator3(10'b1010100011, locator3, alpha34_3_x_locator3);
  gfmult gfm_alpha35_0_x_locator0(10'b0000000001, locator0, alpha35_0_x_locator0);
  gfmult gfm_alpha35_1_x_locator1(10'b1110001011, locator1, alpha35_1_x_locator1);
  gfmult gfm_alpha35_2_x_locator2(10'b1110000111, locator2, alpha35_2_x_locator2);
  gfmult gfm_alpha35_3_x_locator3(10'b0111010111, locator3, alpha35_3_x_locator3);
  gfmult gfm_alpha36_0_x_locator0(10'b0000000001, locator0, alpha36_0_x_locator0);
  gfmult gfm_alpha36_1_x_locator1(10'b1111000001, locator1, alpha36_1_x_locator1);
  gfmult gfm_alpha36_2_x_locator2(10'b1111100111, locator2, alpha36_2_x_locator2);
  gfmult gfm_alpha36_3_x_locator3(10'b1110111101, locator3, alpha36_3_x_locator3);
  gfmult gfm_alpha37_0_x_locator0(10'b0000000001, locator0, alpha37_0_x_locator0);
  gfmult gfm_alpha37_1_x_locator1(10'b1111100100, locator1, alpha37_1_x_locator1);
  gfmult gfm_alpha37_2_x_locator2(10'b1111111111, locator2, alpha37_2_x_locator2);
  gfmult gfm_alpha37_3_x_locator3(10'b1011110010, locator3, alpha37_3_x_locator3);
  gfmult gfm_alpha38_0_x_locator0(10'b0000000001, locator0, alpha38_0_x_locator0);
  gfmult gfm_alpha38_1_x_locator1(10'b0111110010, locator1, alpha38_1_x_locator1);
  gfmult gfm_alpha38_2_x_locator2(10'b1111111001, locator2, alpha38_2_x_locator2);
  gfmult gfm_alpha38_3_x_locator3(10'b0101011100, locator3, alpha38_3_x_locator3);
  gfmult gfm_alpha39_0_x_locator0(10'b0000000001, locator0, alpha39_0_x_locator0);
  gfmult gfm_alpha39_1_x_locator1(10'b0011111001, locator1, alpha39_1_x_locator1);
  gfmult gfm_alpha39_2_x_locator2(10'b0111111100, locator2, alpha39_2_x_locator2);
  gfmult gfm_alpha39_3_x_locator3(10'b1000101111, locator3, alpha39_3_x_locator3);
  gfmult gfm_alpha40_0_x_locator0(10'b0000000001, locator0, alpha40_0_x_locator0);
  gfmult gfm_alpha40_1_x_locator1(10'b1001111000, locator1, alpha40_1_x_locator1);
  gfmult gfm_alpha40_2_x_locator2(10'b0001111111, locator2, alpha40_2_x_locator2);
  gfmult gfm_alpha40_3_x_locator3(10'b1111000010, locator3, alpha40_3_x_locator3);
  gfmult gfm_alpha41_0_x_locator0(10'b0000000001, locator0, alpha41_0_x_locator0);
  gfmult gfm_alpha41_1_x_locator1(10'b0100111100, locator1, alpha41_1_x_locator1);
  gfmult gfm_alpha41_2_x_locator2(10'b1100011001, locator2, alpha41_2_x_locator2);
  gfmult gfm_alpha41_3_x_locator3(10'b0101111010, locator3, alpha41_3_x_locator3);
  gfmult gfm_alpha42_0_x_locator0(10'b0000000001, locator0, alpha42_0_x_locator0);
  gfmult gfm_alpha42_1_x_locator1(10'b0010011110, locator1, alpha42_1_x_locator1);
  gfmult gfm_alpha42_2_x_locator2(10'b0111000100, locator2, alpha42_2_x_locator2);
  gfmult gfm_alpha42_3_x_locator3(10'b0100101101, locator3, alpha42_3_x_locator3);
  gfmult gfm_alpha43_0_x_locator0(10'b0000000001, locator0, alpha43_0_x_locator0);
  gfmult gfm_alpha43_1_x_locator1(10'b0001001111, locator1, alpha43_1_x_locator1);
  gfmult gfm_alpha43_2_x_locator2(10'b0001110001, locator2, alpha43_2_x_locator2);
  gfmult gfm_alpha43_3_x_locator3(10'b1010100000, locator3, alpha43_3_x_locator3);
  gfmult gfm_alpha44_0_x_locator0(10'b0000000001, locator0, alpha44_0_x_locator0);
  gfmult gfm_alpha44_1_x_locator1(10'b1000100011, locator1, alpha44_1_x_locator1);
  gfmult gfm_alpha44_2_x_locator2(10'b0100011110, locator2, alpha44_2_x_locator2);
  gfmult gfm_alpha44_3_x_locator3(10'b0001010100, locator3, alpha44_3_x_locator3);
  gfmult gfm_alpha45_0_x_locator0(10'b0000000001, locator0, alpha45_0_x_locator0);
  gfmult gfm_alpha45_1_x_locator1(10'b1100010101, locator1, alpha45_1_x_locator1);
  gfmult gfm_alpha45_2_x_locator2(10'b1001000011, locator2, alpha45_2_x_locator2);
  gfmult gfm_alpha45_3_x_locator3(10'b1000001110, locator3, alpha45_3_x_locator3);
  gfmult gfm_alpha46_0_x_locator0(10'b0000000001, locator0, alpha46_0_x_locator0);
  gfmult gfm_alpha46_1_x_locator1(10'b1110001110, locator1, alpha46_1_x_locator1);
  gfmult gfm_alpha46_2_x_locator2(10'b1110010110, locator2, alpha46_2_x_locator2);
  gfmult gfm_alpha46_3_x_locator3(10'b1101000111, locator3, alpha46_3_x_locator3);
  gfmult gfm_alpha47_0_x_locator0(10'b0000000001, locator0, alpha47_0_x_locator0);
  gfmult gfm_alpha47_1_x_locator1(10'b0111000111, locator1, alpha47_1_x_locator1);
  gfmult gfm_alpha47_2_x_locator2(10'b1011100001, locator2, alpha47_2_x_locator2);
  gfmult gfm_alpha47_3_x_locator3(10'b1111101111, locator3, alpha47_3_x_locator3);
  gfmult gfm_alpha48_0_x_locator0(10'b0000000001, locator0, alpha48_0_x_locator0);
  gfmult gfm_alpha48_1_x_locator1(10'b1011100111, locator1, alpha48_1_x_locator1);
  gfmult gfm_alpha48_2_x_locator2(10'b0110111010, locator2, alpha48_2_x_locator2);
  gfmult gfm_alpha48_3_x_locator3(10'b1111111010, locator3, alpha48_3_x_locator3);
  gfmult gfm_alpha49_0_x_locator0(10'b0000000001, locator0, alpha49_0_x_locator0);
  gfmult gfm_alpha49_1_x_locator1(10'b1101110111, locator1, alpha49_1_x_locator1);
  gfmult gfm_alpha49_2_x_locator2(10'b1001101010, locator2, alpha49_2_x_locator2);
  gfmult gfm_alpha49_3_x_locator3(10'b0101111101, locator3, alpha49_3_x_locator3);
  gfmult gfm_alpha50_0_x_locator0(10'b0000000001, locator0, alpha50_0_x_locator0);
  gfmult gfm_alpha50_1_x_locator1(10'b1110111111, locator1, alpha50_1_x_locator1);
  gfmult gfm_alpha50_2_x_locator2(10'b1010011110, locator2, alpha50_2_x_locator2);
  gfmult gfm_alpha50_3_x_locator3(10'b1010101010, locator3, alpha50_3_x_locator3);
  gfmult gfm_alpha51_0_x_locator0(10'b0000000001, locator0, alpha51_0_x_locator0);
  gfmult gfm_alpha51_1_x_locator1(10'b1111011011, locator1, alpha51_1_x_locator1);
  gfmult gfm_alpha51_2_x_locator2(10'b1010100011, locator2, alpha51_2_x_locator2);
  gfmult gfm_alpha51_3_x_locator3(10'b0101010111, locator3, alpha51_3_x_locator3);
  gfmult gfm_alpha52_0_x_locator0(10'b0000000001, locator0, alpha52_0_x_locator0);
  gfmult gfm_alpha52_1_x_locator1(10'b1111101001, locator1, alpha52_1_x_locator1);
  gfmult gfm_alpha52_2_x_locator2(10'b1110101110, locator2, alpha52_2_x_locator2);
  gfmult gfm_alpha52_3_x_locator3(10'b1110101101, locator3, alpha52_3_x_locator3);
  gfmult gfm_alpha53_0_x_locator0(10'b0000000001, locator0, alpha53_0_x_locator0);
  gfmult gfm_alpha53_1_x_locator1(10'b1111110000, locator1, alpha53_1_x_locator1);
  gfmult gfm_alpha53_2_x_locator2(10'b1011101111, locator2, alpha53_2_x_locator2);
  gfmult gfm_alpha53_3_x_locator3(10'b1011110000, locator3, alpha53_3_x_locator3);
  gfmult gfm_alpha54_0_x_locator0(10'b0000000001, locator0, alpha54_0_x_locator0);
  gfmult gfm_alpha54_1_x_locator1(10'b0111111000, locator1, alpha54_1_x_locator1);
  gfmult gfm_alpha54_2_x_locator2(10'b1110111101, locator2, alpha54_2_x_locator2);
  gfmult gfm_alpha54_3_x_locator3(10'b0001011110, locator3, alpha54_3_x_locator3);
  gfmult gfm_alpha55_0_x_locator0(10'b0000000001, locator0, alpha55_0_x_locator0);
  gfmult gfm_alpha55_1_x_locator1(10'b0011111100, locator1, alpha55_1_x_locator1);
  gfmult gfm_alpha55_2_x_locator2(10'b0111101101, locator2, alpha55_2_x_locator2);
  gfmult gfm_alpha55_3_x_locator3(10'b1100001101, locator3, alpha55_3_x_locator3);
  gfmult gfm_alpha56_0_x_locator0(10'b0000000001, locator0, alpha56_0_x_locator0);
  gfmult gfm_alpha56_1_x_locator1(10'b0001111110, locator1, alpha56_1_x_locator1);
  gfmult gfm_alpha56_2_x_locator2(10'b0101111001, locator2, alpha56_2_x_locator2);
  gfmult gfm_alpha56_3_x_locator3(10'b1011100100, locator3, alpha56_3_x_locator3);
  gfmult gfm_alpha57_0_x_locator0(10'b0000000001, locator0, alpha57_0_x_locator0);
  gfmult gfm_alpha57_1_x_locator1(10'b0000111111, locator1, alpha57_1_x_locator1);
  gfmult gfm_alpha57_2_x_locator2(10'b0101011100, locator2, alpha57_2_x_locator2);
  gfmult gfm_alpha57_3_x_locator3(10'b1001011000, locator3, alpha57_3_x_locator3);
  gfmult gfm_alpha58_0_x_locator0(10'b0000000001, locator0, alpha58_0_x_locator0);
  gfmult gfm_alpha58_1_x_locator1(10'b1000011011, locator1, alpha58_1_x_locator1);
  gfmult gfm_alpha58_2_x_locator2(10'b0001010111, locator2, alpha58_2_x_locator2);
  gfmult gfm_alpha58_3_x_locator3(10'b0001001011, locator3, alpha58_3_x_locator3);
  gfmult gfm_alpha59_0_x_locator0(10'b0000000001, locator0, alpha59_0_x_locator0);
  gfmult gfm_alpha59_1_x_locator1(10'b1100001001, locator1, alpha59_1_x_locator1);
  gfmult gfm_alpha59_2_x_locator2(10'b1100010011, locator2, alpha59_2_x_locator2);
  gfmult gfm_alpha59_3_x_locator3(10'b0110001010, locator3, alpha59_3_x_locator3);
  gfmult gfm_alpha60_0_x_locator0(10'b0000000001, locator0, alpha60_0_x_locator0);
  gfmult gfm_alpha60_1_x_locator1(10'b1110000000, locator1, alpha60_1_x_locator1);
  gfmult gfm_alpha60_2_x_locator2(10'b1111000010, locator2, alpha60_2_x_locator2);
  gfmult gfm_alpha60_3_x_locator3(10'b0100110011, locator3, alpha60_3_x_locator3);
  gfmult gfm_alpha61_0_x_locator0(10'b0000000001, locator0, alpha61_0_x_locator0);
  gfmult gfm_alpha61_1_x_locator1(10'b0111000000, locator1, alpha61_1_x_locator1);
  gfmult gfm_alpha61_2_x_locator2(10'b1011110100, locator2, alpha61_2_x_locator2);
  gfmult gfm_alpha61_3_x_locator3(10'b0110100101, locator3, alpha61_3_x_locator3);
  gfmult gfm_alpha62_0_x_locator0(10'b0000000001, locator0, alpha62_0_x_locator0);
  gfmult gfm_alpha62_1_x_locator1(10'b0011100000, locator1, alpha62_1_x_locator1);
  gfmult gfm_alpha62_2_x_locator2(10'b0010111101, locator2, alpha62_2_x_locator2);
  gfmult gfm_alpha62_3_x_locator3(10'b1010110001, locator3, alpha62_3_x_locator3);
  gfmult gfm_alpha63_0_x_locator0(10'b0000000001, locator0, alpha63_0_x_locator0);
  gfmult gfm_alpha63_1_x_locator1(10'b0001110000, locator1, alpha63_1_x_locator1);
  gfmult gfm_alpha63_2_x_locator2(10'b0100101101, locator2, alpha63_2_x_locator2);
  gfmult gfm_alpha63_3_x_locator3(10'b0011010111, locator3, alpha63_3_x_locator3);
  gfmult gfm_alpha64_0_x_locator0(10'b0000000001, locator0, alpha64_0_x_locator0);
  gfmult gfm_alpha64_1_x_locator1(10'b0000111000, locator1, alpha64_1_x_locator1);
  gfmult gfm_alpha64_2_x_locator2(10'b0101001001, locator2, alpha64_2_x_locator2);
  gfmult gfm_alpha64_3_x_locator3(10'b1110011101, locator3, alpha64_3_x_locator3);
  gfmult gfm_alpha65_0_x_locator0(10'b0000000001, locator0, alpha65_0_x_locator0);
  gfmult gfm_alpha65_1_x_locator1(10'b0000011100, locator1, alpha65_1_x_locator1);
  gfmult gfm_alpha65_2_x_locator2(10'b0101010000, locator2, alpha65_2_x_locator2);
  gfmult gfm_alpha65_3_x_locator3(10'b1011110110, locator3, alpha65_3_x_locator3);
  gfmult gfm_alpha66_0_x_locator0(10'b0000000001, locator0, alpha66_0_x_locator0);
  gfmult gfm_alpha66_1_x_locator1(10'b0000001110, locator1, alpha66_1_x_locator1);
  gfmult gfm_alpha66_2_x_locator2(10'b0001010100, locator2, alpha66_2_x_locator2);
  gfmult gfm_alpha66_3_x_locator3(10'b1101011000, locator3, alpha66_3_x_locator3);
  gfmult gfm_alpha67_0_x_locator0(10'b0000000001, locator0, alpha67_0_x_locator0);
  gfmult gfm_alpha67_1_x_locator1(10'b0000000111, locator1, alpha67_1_x_locator1);
  gfmult gfm_alpha67_2_x_locator2(10'b0000010101, locator2, alpha67_2_x_locator2);
  gfmult gfm_alpha67_3_x_locator3(10'b0001101011, locator3, alpha67_3_x_locator3);
  gfmult gfm_alpha68_0_x_locator0(10'b0000000001, locator0, alpha68_0_x_locator0);
  gfmult gfm_alpha68_1_x_locator1(10'b1000000111, locator1, alpha68_1_x_locator1);
  gfmult gfm_alpha68_2_x_locator2(10'b0100000111, locator2, alpha68_2_x_locator2);
  gfmult gfm_alpha68_3_x_locator3(10'b0110001110, locator3, alpha68_3_x_locator3);
  gfmult gfm_alpha69_0_x_locator0(10'b0000000001, locator0, alpha69_0_x_locator0);
  gfmult gfm_alpha69_1_x_locator1(10'b1100000111, locator1, alpha69_1_x_locator1);
  gfmult gfm_alpha69_2_x_locator2(10'b1101000111, locator2, alpha69_2_x_locator2);
  gfmult gfm_alpha69_3_x_locator3(10'b1100110111, locator3, alpha69_3_x_locator3);
  gfmult gfm_alpha70_0_x_locator0(10'b0000000001, locator0, alpha70_0_x_locator0);
  gfmult gfm_alpha70_1_x_locator1(10'b1110000111, locator1, alpha70_1_x_locator1);
  gfmult gfm_alpha70_2_x_locator2(10'b1111010111, locator2, alpha70_2_x_locator2);
  gfmult gfm_alpha70_3_x_locator3(10'b1111100001, locator3, alpha70_3_x_locator3);
  gfmult gfm_alpha71_0_x_locator0(10'b0000000001, locator0, alpha71_0_x_locator0);
  gfmult gfm_alpha71_1_x_locator1(10'b1111000111, locator1, alpha71_1_x_locator1);
  gfmult gfm_alpha71_2_x_locator2(10'b1111110011, locator2, alpha71_2_x_locator2);
  gfmult gfm_alpha71_3_x_locator3(10'b0011111101, locator3, alpha71_3_x_locator3);
  gfmult gfm_alpha72_0_x_locator0(10'b0000000001, locator0, alpha72_0_x_locator0);
  gfmult gfm_alpha72_1_x_locator1(10'b1111100111, locator1, alpha72_1_x_locator1);
  gfmult gfm_alpha72_2_x_locator2(10'b1111111010, locator2, alpha72_2_x_locator2);
  gfmult gfm_alpha72_3_x_locator3(10'b1010011010, locator3, alpha72_3_x_locator3);
  gfmult gfm_alpha73_0_x_locator0(10'b0000000001, locator0, alpha73_0_x_locator0);
  gfmult gfm_alpha73_1_x_locator1(10'b1111110111, locator1, alpha73_1_x_locator1);
  gfmult gfm_alpha73_2_x_locator2(10'b1011111010, locator2, alpha73_2_x_locator2);
  gfmult gfm_alpha73_3_x_locator3(10'b0101010001, locator3, alpha73_3_x_locator3);
  gfmult gfm_alpha74_0_x_locator0(10'b0000000001, locator0, alpha74_0_x_locator0);
  gfmult gfm_alpha74_1_x_locator1(10'b1111111111, locator1, alpha74_1_x_locator1);
  gfmult gfm_alpha74_2_x_locator2(10'b1010111010, locator2, alpha74_2_x_locator2);
  gfmult gfm_alpha74_3_x_locator3(10'b0010101011, locator3, alpha74_3_x_locator3);
  gfmult gfm_alpha75_0_x_locator0(10'b0000000001, locator0, alpha75_0_x_locator0);
  gfmult gfm_alpha75_1_x_locator1(10'b1111111011, locator1, alpha75_1_x_locator1);
  gfmult gfm_alpha75_2_x_locator2(10'b1010101010, locator2, alpha75_2_x_locator2);
  gfmult gfm_alpha75_3_x_locator3(10'b0110010110, locator3, alpha75_3_x_locator3);
  gfmult gfm_alpha76_0_x_locator0(10'b0000000001, locator0, alpha76_0_x_locator0);
  gfmult gfm_alpha76_1_x_locator1(10'b1111111001, locator1, alpha76_1_x_locator1);
  gfmult gfm_alpha76_2_x_locator2(10'b1010101110, locator2, alpha76_2_x_locator2);
  gfmult gfm_alpha76_3_x_locator3(10'b1100110100, locator3, alpha76_3_x_locator3);
  gfmult gfm_alpha77_0_x_locator0(10'b0000000001, locator0, alpha77_0_x_locator0);
  gfmult gfm_alpha77_1_x_locator1(10'b1111111000, locator1, alpha77_1_x_locator1);
  gfmult gfm_alpha77_2_x_locator2(10'b1010101111, locator2, alpha77_2_x_locator2);
  gfmult gfm_alpha77_3_x_locator3(10'b1001100010, locator3, alpha77_3_x_locator3);
  gfmult gfm_alpha78_0_x_locator0(10'b0000000001, locator0, alpha78_0_x_locator0);
  gfmult gfm_alpha78_1_x_locator1(10'b0111111100, locator1, alpha78_1_x_locator1);
  gfmult gfm_alpha78_2_x_locator2(10'b1110101101, locator2, alpha78_2_x_locator2);
  gfmult gfm_alpha78_3_x_locator3(10'b0101001110, locator3, alpha78_3_x_locator3);
  gfmult gfm_alpha79_0_x_locator0(10'b0000000001, locator0, alpha79_0_x_locator0);
  gfmult gfm_alpha79_1_x_locator1(10'b0011111110, locator1, alpha79_1_x_locator1);
  gfmult gfm_alpha79_2_x_locator2(10'b0111101001, locator2, alpha79_2_x_locator2);
  gfmult gfm_alpha79_3_x_locator3(10'b1100101111, locator3, alpha79_3_x_locator3);
  gfmult gfm_alpha80_0_x_locator0(10'b0000000001, locator0, alpha80_0_x_locator0);
  gfmult gfm_alpha80_1_x_locator1(10'b0001111111, locator1, alpha80_1_x_locator1);
  gfmult gfm_alpha80_2_x_locator2(10'b0101111000, locator2, alpha80_2_x_locator2);
  gfmult gfm_alpha80_3_x_locator3(10'b1111100010, locator3, alpha80_3_x_locator3);
  gfmult gfm_alpha81_0_x_locator0(10'b0000000001, locator0, alpha81_0_x_locator0);
  gfmult gfm_alpha81_1_x_locator1(10'b1000111011, locator1, alpha81_1_x_locator1);
  gfmult gfm_alpha81_2_x_locator2(10'b0001011110, locator2, alpha81_2_x_locator2);
  gfmult gfm_alpha81_3_x_locator3(10'b0101111110, locator3, alpha81_3_x_locator3);
  gfmult gfm_alpha82_0_x_locator0(10'b0000000001, locator0, alpha82_0_x_locator0);
  gfmult gfm_alpha82_1_x_locator1(10'b1100011001, locator1, alpha82_1_x_locator1);
  gfmult gfm_alpha82_2_x_locator2(10'b1000010011, locator2, alpha82_2_x_locator2);
  gfmult gfm_alpha82_3_x_locator3(10'b1100101001, locator3, alpha82_3_x_locator3);
  gfmult gfm_alpha83_0_x_locator0(10'b0000000001, locator0, alpha83_0_x_locator0);
  gfmult gfm_alpha83_1_x_locator1(10'b1110001000, locator1, alpha83_1_x_locator1);
  gfmult gfm_alpha83_2_x_locator2(10'b1110000010, locator2, alpha83_2_x_locator2);
  gfmult gfm_alpha83_3_x_locator3(10'b0011100100, locator3, alpha83_3_x_locator3);
  gfmult gfm_alpha84_0_x_locator0(10'b0000000001, locator0, alpha84_0_x_locator0);
  gfmult gfm_alpha84_1_x_locator1(10'b0111000100, locator1, alpha84_1_x_locator1);
  gfmult gfm_alpha84_2_x_locator2(10'b1011100100, locator2, alpha84_2_x_locator2);
  gfmult gfm_alpha84_3_x_locator3(10'b1000011000, locator3, alpha84_3_x_locator3);
  gfmult gfm_alpha85_0_x_locator0(10'b0000000001, locator0, alpha85_0_x_locator0);
  gfmult gfm_alpha85_1_x_locator1(10'b0011100010, locator1, alpha85_1_x_locator1);
  gfmult gfm_alpha85_2_x_locator2(10'b0010111001, locator2, alpha85_2_x_locator2);
  gfmult gfm_alpha85_3_x_locator3(10'b0001000011, locator3, alpha85_3_x_locator3);
  gfmult gfm_alpha86_0_x_locator0(10'b0000000001, locator0, alpha86_0_x_locator0);
  gfmult gfm_alpha86_1_x_locator1(10'b0001110001, locator1, alpha86_1_x_locator1);
  gfmult gfm_alpha86_2_x_locator2(10'b0100101100, locator2, alpha86_2_x_locator2);
  gfmult gfm_alpha86_3_x_locator3(10'b0110001011, locator3, alpha86_3_x_locator3);
  gfmult gfm_alpha87_0_x_locator0(10'b0000000001, locator0, alpha87_0_x_locator0);
  gfmult gfm_alpha87_1_x_locator1(10'b1000111100, locator1, alpha87_1_x_locator1);
  gfmult gfm_alpha87_2_x_locator2(10'b0001001011, locator2, alpha87_2_x_locator2);
  gfmult gfm_alpha87_3_x_locator3(10'b0110110010, locator3, alpha87_3_x_locator3);
  gfmult gfm_alpha88_0_x_locator0(10'b0000000001, locator0, alpha88_0_x_locator0);
  gfmult gfm_alpha88_1_x_locator1(10'b0100011110, locator1, alpha88_1_x_locator1);
  gfmult gfm_alpha88_2_x_locator2(10'b1100010100, locator2, alpha88_2_x_locator2);
  gfmult gfm_alpha88_3_x_locator3(10'b0100110100, locator3, alpha88_3_x_locator3);
  gfmult gfm_alpha89_0_x_locator0(10'b0000000001, locator0, alpha89_0_x_locator0);
  gfmult gfm_alpha89_1_x_locator1(10'b0010001111, locator1, alpha89_1_x_locator1);
  gfmult gfm_alpha89_2_x_locator2(10'b0011000101, locator2, alpha89_2_x_locator2);
  gfmult gfm_alpha89_3_x_locator3(10'b1000100010, locator3, alpha89_3_x_locator3);
  gfmult gfm_alpha90_0_x_locator0(10'b0000000001, locator0, alpha90_0_x_locator0);
  gfmult gfm_alpha90_1_x_locator1(10'b1001000011, locator1, alpha90_1_x_locator1);
  gfmult gfm_alpha90_2_x_locator2(10'b0100110011, locator2, alpha90_2_x_locator2);
  gfmult gfm_alpha90_3_x_locator3(10'b0101000110, locator3, alpha90_3_x_locator3);
  gfmult gfm_alpha91_0_x_locator0(10'b0000000001, locator0, alpha91_0_x_locator0);
  gfmult gfm_alpha91_1_x_locator1(10'b1100100101, locator1, alpha91_1_x_locator1);
  gfmult gfm_alpha91_2_x_locator2(10'b1101001010, locator2, alpha91_2_x_locator2);
  gfmult gfm_alpha91_3_x_locator3(10'b1100101110, locator3, alpha91_3_x_locator3);
  gfmult gfm_alpha92_0_x_locator0(10'b0000000001, locator0, alpha92_0_x_locator0);
  gfmult gfm_alpha92_1_x_locator1(10'b1110010110, locator1, alpha92_1_x_locator1);
  gfmult gfm_alpha92_2_x_locator2(10'b1011010110, locator2, alpha92_2_x_locator2);
  gfmult gfm_alpha92_3_x_locator3(10'b1101100011, locator3, alpha92_3_x_locator3);
  gfmult gfm_alpha93_0_x_locator0(10'b0000000001, locator0, alpha93_0_x_locator0);
  gfmult gfm_alpha93_1_x_locator1(10'b0111001011, locator1, alpha93_1_x_locator1);
  gfmult gfm_alpha93_2_x_locator2(10'b1010110001, locator2, alpha93_2_x_locator2);
  gfmult gfm_alpha93_3_x_locator3(10'b0111101111, locator3, alpha93_3_x_locator3);
  gfmult gfm_alpha94_0_x_locator0(10'b0000000001, locator0, alpha94_0_x_locator0);
  gfmult gfm_alpha94_1_x_locator1(10'b1011100001, locator1, alpha94_1_x_locator1);
  gfmult gfm_alpha94_2_x_locator2(10'b0110101110, locator2, alpha94_2_x_locator2);
  gfmult gfm_alpha94_3_x_locator3(10'b1110111010, locator3, alpha94_3_x_locator3);
  gfmult gfm_alpha95_0_x_locator0(10'b0000000001, locator0, alpha95_0_x_locator0);
  gfmult gfm_alpha95_1_x_locator1(10'b1101110100, locator1, alpha95_1_x_locator1);
  gfmult gfm_alpha95_2_x_locator2(10'b1001101111, locator2, alpha95_2_x_locator2);
  gfmult gfm_alpha95_3_x_locator3(10'b0101110101, locator3, alpha95_3_x_locator3);
  gfmult gfm_alpha96_0_x_locator0(10'b0000000001, locator0, alpha96_0_x_locator0);
  gfmult gfm_alpha96_1_x_locator1(10'b0110111010, locator1, alpha96_1_x_locator1);
  gfmult gfm_alpha96_2_x_locator2(10'b1110011101, locator2, alpha96_2_x_locator2);
  gfmult gfm_alpha96_3_x_locator3(10'b1010101011, locator3, alpha96_3_x_locator3);
  gfmult gfm_alpha97_0_x_locator0(10'b0000000001, locator0, alpha97_0_x_locator0);
  gfmult gfm_alpha97_1_x_locator1(10'b0011011101, locator1, alpha97_1_x_locator1);
  gfmult gfm_alpha97_2_x_locator2(10'b0111100101, locator2, alpha97_2_x_locator2);
  gfmult gfm_alpha97_3_x_locator3(10'b0111010110, locator3, alpha97_3_x_locator3);
  gfmult gfm_alpha98_0_x_locator0(10'b0000000001, locator0, alpha98_0_x_locator0);
  gfmult gfm_alpha98_1_x_locator1(10'b1001101010, locator1, alpha98_1_x_locator1);
  gfmult gfm_alpha98_2_x_locator2(10'b0101111011, locator2, alpha98_2_x_locator2);
  gfmult gfm_alpha98_3_x_locator3(10'b1100111100, locator3, alpha98_3_x_locator3);
  gfmult gfm_alpha99_0_x_locator0(10'b0000000001, locator0, alpha99_0_x_locator0);
  gfmult gfm_alpha99_1_x_locator1(10'b0100110101, locator1, alpha99_1_x_locator1);
  gfmult gfm_alpha99_2_x_locator2(10'b1101011000, locator2, alpha99_2_x_locator2);
  gfmult gfm_alpha99_3_x_locator3(10'b1001100011, locator3, alpha99_3_x_locator3);
  gfmult gfm_alpha100_0_x_locator0(10'b0000000001, locator0, alpha100_0_x_locator0);
  gfmult gfm_alpha100_1_x_locator1(10'b1010011110, locator1, alpha100_1_x_locator1);
  gfmult gfm_alpha100_2_x_locator2(10'b0011010110, locator2, alpha100_2_x_locator2);
  gfmult gfm_alpha100_3_x_locator3(10'b0111001111, locator3, alpha100_3_x_locator3);
  gfmult gfm_alpha101_0_x_locator0(10'b0000000001, locator0, alpha101_0_x_locator0);
  gfmult gfm_alpha101_1_x_locator1(10'b0101001111, locator1, alpha101_1_x_locator1);
  gfmult gfm_alpha101_2_x_locator2(10'b1000110001, locator2, alpha101_2_x_locator2);
  gfmult gfm_alpha101_3_x_locator3(10'b1110111110, locator3, alpha101_3_x_locator3);
  gfmult gfm_alpha102_0_x_locator0(10'b0000000001, locator0, alpha102_0_x_locator0);
  gfmult gfm_alpha102_1_x_locator1(10'b1010100011, locator1, alpha102_1_x_locator1);
  gfmult gfm_alpha102_2_x_locator2(10'b0110001110, locator2, alpha102_2_x_locator2);
  gfmult gfm_alpha102_3_x_locator3(10'b1101110001, locator3, alpha102_3_x_locator3);
  gfmult gfm_alpha103_0_x_locator0(10'b0000000001, locator0, alpha103_0_x_locator0);
  gfmult gfm_alpha103_1_x_locator1(10'b1101010101, locator1, alpha103_1_x_locator1);
  gfmult gfm_alpha103_2_x_locator2(10'b1001100111, locator2, alpha103_2_x_locator2);
  gfmult gfm_alpha103_3_x_locator3(10'b0011101111, locator3, alpha103_3_x_locator3);
  gfmult gfm_alpha104_0_x_locator0(10'b0000000001, locator0, alpha104_0_x_locator0);
  gfmult gfm_alpha104_1_x_locator1(10'b1110101110, locator1, alpha104_1_x_locator1);
  gfmult gfm_alpha104_2_x_locator2(10'b1110011111, locator2, alpha104_2_x_locator2);
  gfmult gfm_alpha104_3_x_locator3(10'b1110011010, locator3, alpha104_3_x_locator3);
  gfmult gfm_alpha105_0_x_locator0(10'b0000000001, locator0, alpha105_0_x_locator0);
  gfmult gfm_alpha105_1_x_locator1(10'b0111010111, locator1, alpha105_1_x_locator1);
  gfmult gfm_alpha105_2_x_locator2(10'b1111100001, locator2, alpha105_2_x_locator2);
  gfmult gfm_alpha105_3_x_locator3(10'b0101110001, locator3, alpha105_3_x_locator3);
  gfmult gfm_alpha106_0_x_locator0(10'b0000000001, locator0, alpha106_0_x_locator0);
  gfmult gfm_alpha106_1_x_locator1(10'b1011101111, locator1, alpha106_1_x_locator1);
  gfmult gfm_alpha106_2_x_locator2(10'b0111111010, locator2, alpha106_2_x_locator2);
  gfmult gfm_alpha106_3_x_locator3(10'b0010101111, locator3, alpha106_3_x_locator3);
  gfmult gfm_alpha107_0_x_locator0(10'b0000000001, locator0, alpha107_0_x_locator0);
  gfmult gfm_alpha107_1_x_locator1(10'b1101110011, locator1, alpha107_1_x_locator1);
  gfmult gfm_alpha107_2_x_locator2(10'b1001111010, locator2, alpha107_2_x_locator2);
  gfmult gfm_alpha107_3_x_locator3(10'b1110010010, locator3, alpha107_3_x_locator3);
  gfmult gfm_alpha108_0_x_locator0(10'b0000000001, locator0, alpha108_0_x_locator0);
  gfmult gfm_alpha108_1_x_locator1(10'b1110111101, locator1, alpha108_1_x_locator1);
  gfmult gfm_alpha108_2_x_locator2(10'b1010011010, locator2, alpha108_2_x_locator2);
  gfmult gfm_alpha108_3_x_locator3(10'b0101110000, locator3, alpha108_3_x_locator3);
  gfmult gfm_alpha109_0_x_locator0(10'b0000000001, locator0, alpha109_0_x_locator0);
  gfmult gfm_alpha109_1_x_locator1(10'b1111011010, locator1, alpha109_1_x_locator1);
  gfmult gfm_alpha109_2_x_locator2(10'b1010100010, locator2, alpha109_2_x_locator2);
  gfmult gfm_alpha109_3_x_locator3(10'b0000101110, locator3, alpha109_3_x_locator3);
  gfmult gfm_alpha110_0_x_locator0(10'b0000000001, locator0, alpha110_0_x_locator0);
  gfmult gfm_alpha110_1_x_locator1(10'b0111101101, locator1, alpha110_1_x_locator1);
  gfmult gfm_alpha110_2_x_locator2(10'b1010101100, locator2, alpha110_2_x_locator2);
  gfmult gfm_alpha110_3_x_locator3(10'b1100000011, locator3, alpha110_3_x_locator3);
  gfmult gfm_alpha111_0_x_locator0(10'b0000000001, locator0, alpha111_0_x_locator0);
  gfmult gfm_alpha111_1_x_locator1(10'b1011110010, locator1, alpha111_1_x_locator1);
  gfmult gfm_alpha111_2_x_locator2(10'b0010101011, locator2, alpha111_2_x_locator2);
  gfmult gfm_alpha111_3_x_locator3(10'b0111100011, locator3, alpha111_3_x_locator3);
  gfmult gfm_alpha112_0_x_locator0(10'b0000000001, locator0, alpha112_0_x_locator0);
  gfmult gfm_alpha112_1_x_locator1(10'b0101111001, locator1, alpha112_1_x_locator1);
  gfmult gfm_alpha112_2_x_locator2(10'b1100101100, locator2, alpha112_2_x_locator2);
  gfmult gfm_alpha112_3_x_locator3(10'b0110111111, locator3, alpha112_3_x_locator3);
  gfmult gfm_alpha113_0_x_locator0(10'b0000000001, locator0, alpha113_0_x_locator0);
  gfmult gfm_alpha113_1_x_locator1(10'b1010111000, locator1, alpha113_1_x_locator1);
  gfmult gfm_alpha113_2_x_locator2(10'b0011001011, locator2, alpha113_2_x_locator2);
  gfmult gfm_alpha113_3_x_locator3(10'b1110110000, locator3, alpha113_3_x_locator3);
  gfmult gfm_alpha114_0_x_locator0(10'b0000000001, locator0, alpha114_0_x_locator0);
  gfmult gfm_alpha114_1_x_locator1(10'b0101011100, locator1, alpha114_1_x_locator1);
  gfmult gfm_alpha114_2_x_locator2(10'b1100110100, locator2, alpha114_2_x_locator2);
  gfmult gfm_alpha114_3_x_locator3(10'b0001110110, locator3, alpha114_3_x_locator3);
  gfmult gfm_alpha115_0_x_locator0(10'b0000000001, locator0, alpha115_0_x_locator0);
  gfmult gfm_alpha115_1_x_locator1(10'b0010101110, locator1, alpha115_1_x_locator1);
  gfmult gfm_alpha115_2_x_locator2(10'b0011001101, locator2, alpha115_2_x_locator2);
  gfmult gfm_alpha115_3_x_locator3(10'b1100001000, locator3, alpha115_3_x_locator3);
  gfmult gfm_alpha116_0_x_locator0(10'b0000000001, locator0, alpha116_0_x_locator0);
  gfmult gfm_alpha116_1_x_locator1(10'b0001010111, locator1, alpha116_1_x_locator1);
  gfmult gfm_alpha116_2_x_locator2(10'b0100110001, locator2, alpha116_2_x_locator2);
  gfmult gfm_alpha116_3_x_locator3(10'b0001100001, locator3, alpha116_3_x_locator3);
  gfmult gfm_alpha117_0_x_locator0(10'b0000000001, locator0, alpha117_0_x_locator0);
  gfmult gfm_alpha117_1_x_locator1(10'b1000101111, locator1, alpha117_1_x_locator1);
  gfmult gfm_alpha117_2_x_locator2(10'b0101001110, locator2, alpha117_2_x_locator2);
  gfmult gfm_alpha117_3_x_locator3(10'b0010001101, locator3, alpha117_3_x_locator3);
  gfmult gfm_alpha118_0_x_locator0(10'b0000000001, locator0, alpha118_0_x_locator0);
  gfmult gfm_alpha118_1_x_locator1(10'b1100010011, locator1, alpha118_1_x_locator1);
  gfmult gfm_alpha118_2_x_locator2(10'b1001010111, locator2, alpha118_2_x_locator2);
  gfmult gfm_alpha118_3_x_locator3(10'b1010010100, locator3, alpha118_3_x_locator3);
  gfmult gfm_alpha119_0_x_locator0(10'b0000000001, locator0, alpha119_0_x_locator0);
  gfmult gfm_alpha119_1_x_locator1(10'b1110001101, locator1, alpha119_1_x_locator1);
  gfmult gfm_alpha119_2_x_locator2(10'b1110010011, locator2, alpha119_2_x_locator2);
  gfmult gfm_alpha119_3_x_locator3(10'b1001010110, locator3, alpha119_3_x_locator3);
  gfmult gfm_alpha120_0_x_locator0(10'b0000000001, locator0, alpha120_0_x_locator0);
  gfmult gfm_alpha120_1_x_locator1(10'b1111000010, locator1, alpha120_1_x_locator1);
  gfmult gfm_alpha120_2_x_locator2(10'b1111100010, locator2, alpha120_2_x_locator2);
  gfmult gfm_alpha120_3_x_locator3(10'b1101001100, locator3, alpha120_3_x_locator3);
  gfmult gfm_alpha121_0_x_locator0(10'b0000000001, locator0, alpha121_0_x_locator0);
  gfmult gfm_alpha121_1_x_locator1(10'b0111100001, locator1, alpha121_1_x_locator1);
  gfmult gfm_alpha121_2_x_locator2(10'b1011111100, locator2, alpha121_2_x_locator2);
  gfmult gfm_alpha121_3_x_locator3(10'b1001101101, locator3, alpha121_3_x_locator3);
  gfmult gfm_alpha122_0_x_locator0(10'b0000000001, locator0, alpha122_0_x_locator0);
  gfmult gfm_alpha122_1_x_locator1(10'b1011110100, locator1, alpha122_1_x_locator1);
  gfmult gfm_alpha122_2_x_locator2(10'b0010111111, locator2, alpha122_2_x_locator2);
  gfmult gfm_alpha122_3_x_locator3(10'b1011001000, locator3, alpha122_3_x_locator3);
  gfmult gfm_alpha123_0_x_locator0(10'b0000000001, locator0, alpha123_0_x_locator0);
  gfmult gfm_alpha123_1_x_locator1(10'b0101111010, locator1, alpha123_1_x_locator1);
  gfmult gfm_alpha123_2_x_locator2(10'b1100101001, locator2, alpha123_2_x_locator2);
  gfmult gfm_alpha123_3_x_locator3(10'b0001011001, locator3, alpha123_3_x_locator3);
  gfmult gfm_alpha124_0_x_locator0(10'b0000000001, locator0, alpha124_0_x_locator0);
  gfmult gfm_alpha124_1_x_locator1(10'b0010111101, locator1, alpha124_1_x_locator1);
  gfmult gfm_alpha124_2_x_locator2(10'b0111001000, locator2, alpha124_2_x_locator2);
  gfmult gfm_alpha124_3_x_locator3(10'b0010001010, locator3, alpha124_3_x_locator3);
  gfmult gfm_alpha125_0_x_locator0(10'b0000000001, locator0, alpha125_0_x_locator0);
  gfmult gfm_alpha125_1_x_locator1(10'b1001011010, locator1, alpha125_1_x_locator1);
  gfmult gfm_alpha125_2_x_locator2(10'b0001110010, locator2, alpha125_2_x_locator2);
  gfmult gfm_alpha125_3_x_locator3(10'b0100010011, locator3, alpha125_3_x_locator3);
  gfmult gfm_alpha126_0_x_locator0(10'b0000000001, locator0, alpha126_0_x_locator0);
  gfmult gfm_alpha126_1_x_locator1(10'b0100101101, locator1, alpha126_1_x_locator1);
  gfmult gfm_alpha126_2_x_locator2(10'b1000011000, locator2, alpha126_2_x_locator2);
  gfmult gfm_alpha126_3_x_locator3(10'b0110100001, locator3, alpha126_3_x_locator3);
  gfmult gfm_alpha127_0_x_locator0(10'b0000000001, locator0, alpha127_0_x_locator0);
  gfmult gfm_alpha127_1_x_locator1(10'b1010010010, locator1, alpha127_1_x_locator1);
  gfmult gfm_alpha127_2_x_locator2(10'b0010000110, locator2, alpha127_2_x_locator2);
  gfmult gfm_alpha127_3_x_locator3(10'b0010110101, locator3, alpha127_3_x_locator3);
  gfmult gfm_alpha128_0_x_locator0(10'b0000000001, locator0, alpha128_0_x_locator0);
  gfmult gfm_alpha128_1_x_locator1(10'b0101001001, locator1, alpha128_1_x_locator1);
  gfmult gfm_alpha128_2_x_locator2(10'b1000100101, locator2, alpha128_2_x_locator2);
  gfmult gfm_alpha128_3_x_locator3(10'b1010010011, locator3, alpha128_3_x_locator3);
  gfmult gfm_alpha129_0_x_locator0(10'b0000000001, locator0, alpha129_0_x_locator0);
  gfmult gfm_alpha129_1_x_locator1(10'b1010100000, locator1, alpha129_1_x_locator1);
  gfmult gfm_alpha129_2_x_locator2(10'b0110001011, locator2, alpha129_2_x_locator2);
  gfmult gfm_alpha129_3_x_locator3(10'b0111010001, locator3, alpha129_3_x_locator3);
  gfmult gfm_alpha130_0_x_locator0(10'b0000000001, locator0, alpha130_0_x_locator0);
  gfmult gfm_alpha130_1_x_locator1(10'b0101010000, locator1, alpha130_1_x_locator1);
  gfmult gfm_alpha130_2_x_locator2(10'b1101100100, locator2, alpha130_2_x_locator2);
  gfmult gfm_alpha130_3_x_locator3(10'b0010111011, locator3, alpha130_3_x_locator3);
  gfmult gfm_alpha131_0_x_locator0(10'b0000000001, locator0, alpha131_0_x_locator0);
  gfmult gfm_alpha131_1_x_locator1(10'b0010101000, locator1, alpha131_1_x_locator1);
  gfmult gfm_alpha131_2_x_locator2(10'b0011011001, locator2, alpha131_2_x_locator2);
  gfmult gfm_alpha131_3_x_locator3(10'b0110010100, locator3, alpha131_3_x_locator3);
  gfmult gfm_alpha132_0_x_locator0(10'b0000000001, locator0, alpha132_0_x_locator0);
  gfmult gfm_alpha132_1_x_locator1(10'b0001010100, locator1, alpha132_1_x_locator1);
  gfmult gfm_alpha132_2_x_locator2(10'b0100110100, locator2, alpha132_2_x_locator2);
  gfmult gfm_alpha132_3_x_locator3(10'b1000110110, locator3, alpha132_3_x_locator3);
  gfmult gfm_alpha133_0_x_locator0(10'b0000000001, locator0, alpha133_0_x_locator0);
  gfmult gfm_alpha133_1_x_locator1(10'b0000101010, locator1, alpha133_1_x_locator1);
  gfmult gfm_alpha133_2_x_locator2(10'b0001001101, locator2, alpha133_2_x_locator2);
  gfmult gfm_alpha133_3_x_locator3(10'b1101000000, locator3, alpha133_3_x_locator3);
  gfmult gfm_alpha134_0_x_locator0(10'b0000000001, locator0, alpha134_0_x_locator0);
  gfmult gfm_alpha134_1_x_locator1(10'b0000010101, locator1, alpha134_1_x_locator1);
  gfmult gfm_alpha134_2_x_locator2(10'b0100010001, locator2, alpha134_2_x_locator2);
  gfmult gfm_alpha134_3_x_locator3(10'b0001101000, locator3, alpha134_3_x_locator3);
  gfmult gfm_alpha135_0_x_locator0(10'b0000000001, locator0, alpha135_0_x_locator0);
  gfmult gfm_alpha135_1_x_locator1(10'b1000001110, locator1, alpha135_1_x_locator1);
  gfmult gfm_alpha135_2_x_locator2(10'b0101000110, locator2, alpha135_2_x_locator2);
  gfmult gfm_alpha135_3_x_locator3(10'b0000001101, locator3, alpha135_3_x_locator3);
  gfmult gfm_alpha136_0_x_locator0(10'b0000000001, locator0, alpha136_0_x_locator0);
  gfmult gfm_alpha136_1_x_locator1(10'b0100000111, locator1, alpha136_1_x_locator1);
  gfmult gfm_alpha136_2_x_locator2(10'b1001010101, locator2, alpha136_2_x_locator2);
  gfmult gfm_alpha136_3_x_locator3(10'b1010000100, locator3, alpha136_3_x_locator3);
  gfmult gfm_alpha137_0_x_locator0(10'b0000000001, locator0, alpha137_0_x_locator0);
  gfmult gfm_alpha137_1_x_locator1(10'b1010000111, locator1, alpha137_1_x_locator1);
  gfmult gfm_alpha137_2_x_locator2(10'b0110010111, locator2, alpha137_2_x_locator2);
  gfmult gfm_alpha137_3_x_locator3(10'b1001010100, locator3, alpha137_3_x_locator3);
  gfmult gfm_alpha138_0_x_locator0(10'b0000000001, locator0, alpha138_0_x_locator0);
  gfmult gfm_alpha138_1_x_locator1(10'b1101000111, locator1, alpha138_1_x_locator1);
  gfmult gfm_alpha138_2_x_locator2(10'b1101100011, locator2, alpha138_2_x_locator2);
  gfmult gfm_alpha138_3_x_locator3(10'b1001001110, locator3, alpha138_3_x_locator3);
  gfmult gfm_alpha139_0_x_locator0(10'b0000000001, locator0, alpha139_0_x_locator0);
  gfmult gfm_alpha139_1_x_locator1(10'b1110100111, locator1, alpha139_1_x_locator1);
  gfmult gfm_alpha139_2_x_locator2(10'b1111011110, locator2, alpha139_2_x_locator2);
  gfmult gfm_alpha139_3_x_locator3(10'b1101001111, locator3, alpha139_3_x_locator3);
  gfmult gfm_alpha140_0_x_locator0(10'b0000000001, locator0, alpha140_0_x_locator0);
  gfmult gfm_alpha140_1_x_locator1(10'b1111010111, locator1, alpha140_1_x_locator1);
  gfmult gfm_alpha140_2_x_locator2(10'b1011110011, locator2, alpha140_2_x_locator2);
  gfmult gfm_alpha140_3_x_locator3(10'b1111101110, locator3, alpha140_3_x_locator3);
  gfmult gfm_alpha141_0_x_locator0(10'b0000000001, locator0, alpha141_0_x_locator0);
  gfmult gfm_alpha141_1_x_locator1(10'b1111101111, locator1, alpha141_1_x_locator1);
  gfmult gfm_alpha141_2_x_locator2(10'b1110111010, locator2, alpha141_2_x_locator2);
  gfmult gfm_alpha141_3_x_locator3(10'b1101111011, locator3, alpha141_3_x_locator3);
  gfmult gfm_alpha142_0_x_locator0(10'b0000000001, locator0, alpha142_0_x_locator0);
  gfmult gfm_alpha142_1_x_locator1(10'b1111110011, locator1, alpha142_1_x_locator1);
  gfmult gfm_alpha142_2_x_locator2(10'b1011101010, locator2, alpha142_2_x_locator2);
  gfmult gfm_alpha142_3_x_locator3(10'b0111101100, locator3, alpha142_3_x_locator3);
  gfmult gfm_alpha143_0_x_locator0(10'b0000000001, locator0, alpha143_0_x_locator0);
  gfmult gfm_alpha143_1_x_locator1(10'b1111111101, locator1, alpha143_1_x_locator1);
  gfmult gfm_alpha143_2_x_locator2(10'b1010111110, locator2, alpha143_2_x_locator2);
  gfmult gfm_alpha143_3_x_locator3(10'b1000111001, locator3, alpha143_3_x_locator3);
  gfmult gfm_alpha144_0_x_locator0(10'b0000000001, locator0, alpha144_0_x_locator0);
  gfmult gfm_alpha144_1_x_locator1(10'b1111111010, locator1, alpha144_1_x_locator1);
  gfmult gfm_alpha144_2_x_locator2(10'b1010101011, locator2, alpha144_2_x_locator2);
  gfmult gfm_alpha144_3_x_locator3(10'b0011000110, locator3, alpha144_3_x_locator3);
  gfmult gfm_alpha145_0_x_locator0(10'b0000000001, locator0, alpha145_0_x_locator0);
  gfmult gfm_alpha145_1_x_locator1(10'b0111111101, locator1, alpha145_1_x_locator1);
  gfmult gfm_alpha145_2_x_locator2(10'b1110101100, locator2, alpha145_2_x_locator2);
  gfmult gfm_alpha145_3_x_locator3(10'b1100011110, locator3, alpha145_3_x_locator3);
  gfmult gfm_alpha146_0_x_locator0(10'b0000000001, locator0, alpha146_0_x_locator0);
  gfmult gfm_alpha146_1_x_locator1(10'b1011111010, locator1, alpha146_1_x_locator1);
  gfmult gfm_alpha146_2_x_locator2(10'b0011101011, locator2, alpha146_2_x_locator2);
  gfmult gfm_alpha146_3_x_locator3(10'b1101100101, locator3, alpha146_3_x_locator3);
  gfmult gfm_alpha147_0_x_locator0(10'b0000000001, locator0, alpha147_0_x_locator0);
  gfmult gfm_alpha147_1_x_locator1(10'b0101111101, locator1, alpha147_1_x_locator1);
  gfmult gfm_alpha147_2_x_locator2(10'b1100111100, locator2, alpha147_2_x_locator2);
  gfmult gfm_alpha147_3_x_locator3(10'b1011101001, locator3, alpha147_3_x_locator3);
  gfmult gfm_alpha148_0_x_locator0(10'b0000000001, locator0, alpha148_0_x_locator0);
  gfmult gfm_alpha148_1_x_locator1(10'b1010111010, locator1, alpha148_1_x_locator1);
  gfmult gfm_alpha148_2_x_locator2(10'b0011001111, locator2, alpha148_2_x_locator2);
  gfmult gfm_alpha148_3_x_locator3(10'b0011011100, locator3, alpha148_3_x_locator3);
  gfmult gfm_alpha149_0_x_locator0(10'b0000000001, locator0, alpha149_0_x_locator0);
  gfmult gfm_alpha149_1_x_locator1(10'b0101011101, locator1, alpha149_1_x_locator1);
  gfmult gfm_alpha149_2_x_locator2(10'b1100110101, locator2, alpha149_2_x_locator2);
  gfmult gfm_alpha149_3_x_locator3(10'b1000011111, locator3, alpha149_3_x_locator3);
  gfmult gfm_alpha150_0_x_locator0(10'b0000000001, locator0, alpha150_0_x_locator0);
  gfmult gfm_alpha150_1_x_locator1(10'b1010101010, locator1, alpha150_1_x_locator1);
  gfmult gfm_alpha150_2_x_locator2(10'b0111001111, locator2, alpha150_2_x_locator2);
  gfmult gfm_alpha150_3_x_locator3(10'b1111000100, locator3, alpha150_3_x_locator3);
  gfmult gfm_alpha151_0_x_locator0(10'b0000000001, locator0, alpha151_0_x_locator0);
  gfmult gfm_alpha151_1_x_locator1(10'b0101010101, locator1, alpha151_1_x_locator1);
  gfmult gfm_alpha151_2_x_locator2(10'b1101110101, locator2, alpha151_2_x_locator2);
  gfmult gfm_alpha151_3_x_locator3(10'b1001111100, locator3, alpha151_3_x_locator3);
  gfmult gfm_alpha152_0_x_locator0(10'b0000000001, locator0, alpha152_0_x_locator0);
  gfmult gfm_alpha152_1_x_locator1(10'b1010101110, locator1, alpha152_1_x_locator1);
  gfmult gfm_alpha152_2_x_locator2(10'b0111011111, locator2, alpha152_2_x_locator2);
  gfmult gfm_alpha152_3_x_locator3(10'b1001001011, locator3, alpha152_3_x_locator3);
  gfmult gfm_alpha153_0_x_locator0(10'b0000000001, locator0, alpha153_0_x_locator0);
  gfmult gfm_alpha153_1_x_locator1(10'b0101010111, locator1, alpha153_1_x_locator1);
  gfmult gfm_alpha153_2_x_locator2(10'b1101110001, locator2, alpha153_2_x_locator2);
  gfmult gfm_alpha153_3_x_locator3(10'b0111001010, locator3, alpha153_3_x_locator3);
  gfmult gfm_alpha154_0_x_locator0(10'b0000000001, locator0, alpha154_0_x_locator0);
  gfmult gfm_alpha154_1_x_locator1(10'b1010101111, locator1, alpha154_1_x_locator1);
  gfmult gfm_alpha154_2_x_locator2(10'b0111011110, locator2, alpha154_2_x_locator2);
  gfmult gfm_alpha154_3_x_locator3(10'b0100111011, locator3, alpha154_3_x_locator3);
  gfmult gfm_alpha155_0_x_locator0(10'b0000000001, locator0, alpha155_0_x_locator0);
  gfmult gfm_alpha155_1_x_locator1(10'b1101010011, locator1, alpha155_1_x_locator1);
  gfmult gfm_alpha155_2_x_locator2(10'b1001110011, locator2, alpha155_2_x_locator2);
  gfmult gfm_alpha155_3_x_locator3(10'b0110100100, locator3, alpha155_3_x_locator3);
  gfmult gfm_alpha156_0_x_locator0(10'b0000000001, locator0, alpha156_0_x_locator0);
  gfmult gfm_alpha156_1_x_locator1(10'b1110101101, locator1, alpha156_1_x_locator1);
  gfmult gfm_alpha156_2_x_locator2(10'b1110011010, locator2, alpha156_2_x_locator2);
  gfmult gfm_alpha156_3_x_locator3(10'b1000110000, locator3, alpha156_3_x_locator3);
  gfmult gfm_alpha157_0_x_locator0(10'b0000000001, locator0, alpha157_0_x_locator0);
  gfmult gfm_alpha157_1_x_locator1(10'b1111010010, locator1, alpha157_1_x_locator1);
  gfmult gfm_alpha157_2_x_locator2(10'b1011100010, locator2, alpha157_2_x_locator2);
  gfmult gfm_alpha157_3_x_locator3(10'b0001000110, locator3, alpha157_3_x_locator3);
  gfmult gfm_alpha158_0_x_locator0(10'b0000000001, locator0, alpha158_0_x_locator0);
  gfmult gfm_alpha158_1_x_locator1(10'b0111101001, locator1, alpha158_1_x_locator1);
  gfmult gfm_alpha158_2_x_locator2(10'b1010111100, locator2, alpha158_2_x_locator2);
  gfmult gfm_alpha158_3_x_locator3(10'b1100001110, locator3, alpha158_3_x_locator3);
  gfmult gfm_alpha159_0_x_locator0(10'b0000000001, locator0, alpha159_0_x_locator0);
  gfmult gfm_alpha159_1_x_locator1(10'b1011110000, locator1, alpha159_1_x_locator1);
  gfmult gfm_alpha159_2_x_locator2(10'b0010101111, locator2, alpha159_2_x_locator2);
  gfmult gfm_alpha159_3_x_locator3(10'b1101100111, locator3, alpha159_3_x_locator3);
  gfmult gfm_alpha160_0_x_locator0(10'b0000000001, locator0, alpha160_0_x_locator0);
  gfmult gfm_alpha160_1_x_locator1(10'b0101111000, locator1, alpha160_1_x_locator1);
  gfmult gfm_alpha160_2_x_locator2(10'b1100101101, locator2, alpha160_2_x_locator2);
  gfmult gfm_alpha160_3_x_locator3(10'b1111101011, locator3, alpha160_3_x_locator3);
  gfmult gfm_alpha161_0_x_locator0(10'b0000000001, locator0, alpha161_0_x_locator0);
  gfmult gfm_alpha161_1_x_locator1(10'b0010111100, locator1, alpha161_1_x_locator1);
  gfmult gfm_alpha161_2_x_locator2(10'b0111001001, locator2, alpha161_2_x_locator2);
  gfmult gfm_alpha161_3_x_locator3(10'b0111111110, locator3, alpha161_3_x_locator3);
  gfmult gfm_alpha162_0_x_locator0(10'b0000000001, locator0, alpha162_0_x_locator0);
  gfmult gfm_alpha162_1_x_locator1(10'b0001011110, locator1, alpha162_1_x_locator1);
  gfmult gfm_alpha162_2_x_locator2(10'b0101110000, locator2, alpha162_2_x_locator2);
  gfmult gfm_alpha162_3_x_locator3(10'b1100111001, locator3, alpha162_3_x_locator3);
  gfmult gfm_alpha163_0_x_locator0(10'b0000000001, locator0, alpha163_0_x_locator0);
  gfmult gfm_alpha163_1_x_locator1(10'b0000101111, locator1, alpha163_1_x_locator1);
  gfmult gfm_alpha163_2_x_locator2(10'b0001011100, locator2, alpha163_2_x_locator2);
  gfmult gfm_alpha163_3_x_locator3(10'b0011100110, locator3, alpha163_3_x_locator3);
  gfmult gfm_alpha164_0_x_locator0(10'b0000000001, locator0, alpha164_0_x_locator0);
  gfmult gfm_alpha164_1_x_locator1(10'b1000010011, locator1, alpha164_1_x_locator1);
  gfmult gfm_alpha164_2_x_locator2(10'b0000010111, locator2, alpha164_2_x_locator2);
  gfmult gfm_alpha164_3_x_locator3(10'b1100011010, locator3, alpha164_3_x_locator3);
  gfmult gfm_alpha165_0_x_locator0(10'b0000000001, locator0, alpha165_0_x_locator0);
  gfmult gfm_alpha165_1_x_locator1(10'b1100001101, locator1, alpha165_1_x_locator1);
  gfmult gfm_alpha165_2_x_locator2(10'b1100000011, locator2, alpha165_2_x_locator2);
  gfmult gfm_alpha165_3_x_locator3(10'b0101100001, locator3, alpha165_3_x_locator3);
  gfmult gfm_alpha166_0_x_locator0(10'b0000000001, locator0, alpha166_0_x_locator0);
  gfmult gfm_alpha166_1_x_locator1(10'b1110000010, locator1, alpha166_1_x_locator1);
  gfmult gfm_alpha166_2_x_locator2(10'b1111000110, locator2, alpha166_2_x_locator2);
  gfmult gfm_alpha166_3_x_locator3(10'b0010101101, locator3, alpha166_3_x_locator3);
  gfmult gfm_alpha167_0_x_locator0(10'b0000000001, locator0, alpha167_0_x_locator0);
  gfmult gfm_alpha167_1_x_locator1(10'b0111000001, locator1, alpha167_1_x_locator1);
  gfmult gfm_alpha167_2_x_locator2(10'b1011110101, locator2, alpha167_2_x_locator2);
  gfmult gfm_alpha167_3_x_locator3(10'b1010010000, locator3, alpha167_3_x_locator3);
  gfmult gfm_alpha168_0_x_locator0(10'b0000000001, locator0, alpha168_0_x_locator0);
  gfmult gfm_alpha168_1_x_locator1(10'b1011100100, locator1, alpha168_1_x_locator1);
  gfmult gfm_alpha168_2_x_locator2(10'b0110111111, locator2, alpha168_2_x_locator2);
  gfmult gfm_alpha168_3_x_locator3(10'b0001010010, locator3, alpha168_3_x_locator3);
  gfmult gfm_alpha169_0_x_locator0(10'b0000000001, locator0, alpha169_0_x_locator0);
  gfmult gfm_alpha169_1_x_locator1(10'b0101110010, locator1, alpha169_1_x_locator1);
  gfmult gfm_alpha169_2_x_locator2(10'b1101101001, locator2, alpha169_2_x_locator2);
  gfmult gfm_alpha169_3_x_locator3(10'b0100001000, locator3, alpha169_3_x_locator3);
  gfmult gfm_alpha170_0_x_locator0(10'b0000000001, locator0, alpha170_0_x_locator0);
  gfmult gfm_alpha170_1_x_locator1(10'b0010111001, locator1, alpha170_1_x_locator1);
  gfmult gfm_alpha170_2_x_locator2(10'b0111011000, locator2, alpha170_2_x_locator2);
  gfmult gfm_alpha170_3_x_locator3(10'b0000100001, locator3, alpha170_3_x_locator3);
  gfmult gfm_alpha171_0_x_locator0(10'b0000000001, locator0, alpha171_0_x_locator0);
  gfmult gfm_alpha171_1_x_locator1(10'b1001011000, locator1, alpha171_1_x_locator1);
  gfmult gfm_alpha171_2_x_locator2(10'b0001110110, locator2, alpha171_2_x_locator2);
  gfmult gfm_alpha171_3_x_locator3(10'b0010000101, locator3, alpha171_3_x_locator3);
  gfmult gfm_alpha172_0_x_locator0(10'b0000000001, locator0, alpha172_0_x_locator0);
  gfmult gfm_alpha172_1_x_locator1(10'b0100101100, locator1, alpha172_1_x_locator1);
  gfmult gfm_alpha172_2_x_locator2(10'b1000011001, locator2, alpha172_2_x_locator2);
  gfmult gfm_alpha172_3_x_locator3(10'b1010010101, locator3, alpha172_3_x_locator3);
  gfmult gfm_alpha173_0_x_locator0(10'b0000000001, locator0, alpha173_0_x_locator0);
  gfmult gfm_alpha173_1_x_locator1(10'b0010010110, locator1, alpha173_1_x_locator1);
  gfmult gfm_alpha173_2_x_locator2(10'b0110000100, locator2, alpha173_2_x_locator2);
  gfmult gfm_alpha173_3_x_locator3(10'b1011010111, locator3, alpha173_3_x_locator3);
  gfmult gfm_alpha174_0_x_locator0(10'b0000000001, locator0, alpha174_0_x_locator0);
  gfmult gfm_alpha174_1_x_locator1(10'b0001001011, locator1, alpha174_1_x_locator1);
  gfmult gfm_alpha174_2_x_locator2(10'b0001100001, locator2, alpha174_2_x_locator2);
  gfmult gfm_alpha174_3_x_locator3(10'b1111011101, locator3, alpha174_3_x_locator3);
  gfmult gfm_alpha175_0_x_locator0(10'b0000000001, locator0, alpha175_0_x_locator0);
  gfmult gfm_alpha175_1_x_locator1(10'b1000100001, locator1, alpha175_1_x_locator1);
  gfmult gfm_alpha175_2_x_locator2(10'b0100011010, locator2, alpha175_2_x_locator2);
  gfmult gfm_alpha175_3_x_locator3(10'b1011111110, locator3, alpha175_3_x_locator3);
  gfmult gfm_alpha176_0_x_locator0(10'b0000000001, locator0, alpha176_0_x_locator0);
  gfmult gfm_alpha176_1_x_locator1(10'b1100010100, locator1, alpha176_1_x_locator1);
  gfmult gfm_alpha176_2_x_locator2(10'b1001000010, locator2, alpha176_2_x_locator2);
  gfmult gfm_alpha176_3_x_locator3(10'b1101011001, locator3, alpha176_3_x_locator3);
  gfmult gfm_alpha177_0_x_locator0(10'b0000000001, locator0, alpha177_0_x_locator0);
  gfmult gfm_alpha177_1_x_locator1(10'b0110001010, locator1, alpha177_1_x_locator1);
  gfmult gfm_alpha177_2_x_locator2(10'b1010010100, locator2, alpha177_2_x_locator2);
  gfmult gfm_alpha177_3_x_locator3(10'b0011101010, locator3, alpha177_3_x_locator3);
  gfmult gfm_alpha178_0_x_locator0(10'b0000000001, locator0, alpha178_0_x_locator0);
  gfmult gfm_alpha178_1_x_locator1(10'b0011000101, locator1, alpha178_1_x_locator1);
  gfmult gfm_alpha178_2_x_locator2(10'b0010100101, locator2, alpha178_2_x_locator2);
  gfmult gfm_alpha178_3_x_locator3(10'b0100011111, locator3, alpha178_3_x_locator3);
  gfmult gfm_alpha179_0_x_locator0(10'b0000000001, locator0, alpha179_0_x_locator0);
  gfmult gfm_alpha179_1_x_locator1(10'b1001100110, locator1, alpha179_1_x_locator1);
  gfmult gfm_alpha179_2_x_locator2(10'b0100101011, locator2, alpha179_2_x_locator2);
  gfmult gfm_alpha179_3_x_locator3(10'b1110100100, locator3, alpha179_3_x_locator3);
  gfmult gfm_alpha180_0_x_locator0(10'b0000000001, locator0, alpha180_0_x_locator0);
  gfmult gfm_alpha180_1_x_locator1(10'b0100110011, locator1, alpha180_1_x_locator1);
  gfmult gfm_alpha180_2_x_locator2(10'b1101001100, locator2, alpha180_2_x_locator2);
  gfmult gfm_alpha180_3_x_locator3(10'b1001110000, locator3, alpha180_3_x_locator3);
  gfmult gfm_alpha181_0_x_locator0(10'b0000000001, locator0, alpha181_0_x_locator0);
  gfmult gfm_alpha181_1_x_locator1(10'b1010011101, locator1, alpha181_1_x_locator1);
  gfmult gfm_alpha181_2_x_locator2(10'b0011010011, locator2, alpha181_2_x_locator2);
  gfmult gfm_alpha181_3_x_locator3(10'b0001001110, locator3, alpha181_3_x_locator3);
  gfmult gfm_alpha182_0_x_locator0(10'b0000000001, locator0, alpha182_0_x_locator0);
  gfmult gfm_alpha182_1_x_locator1(10'b1101001010, locator1, alpha182_1_x_locator1);
  gfmult gfm_alpha182_2_x_locator2(10'b1100110010, locator2, alpha182_2_x_locator2);
  gfmult gfm_alpha182_3_x_locator3(10'b1100001111, locator3, alpha182_3_x_locator3);
  gfmult gfm_alpha183_0_x_locator0(10'b0000000001, locator0, alpha183_0_x_locator0);
  gfmult gfm_alpha183_1_x_locator1(10'b0110100101, locator1, alpha183_1_x_locator1);
  gfmult gfm_alpha183_2_x_locator2(10'b1011001000, locator2, alpha183_2_x_locator2);
  gfmult gfm_alpha183_3_x_locator3(10'b1111100110, locator3, alpha183_3_x_locator3);
  gfmult gfm_alpha184_0_x_locator0(10'b0000000001, locator0, alpha184_0_x_locator0);
  gfmult gfm_alpha184_1_x_locator1(10'b1011010110, locator1, alpha184_1_x_locator1);
  gfmult gfm_alpha184_2_x_locator2(10'b0010110010, locator2, alpha184_2_x_locator2);
  gfmult gfm_alpha184_3_x_locator3(10'b1101111010, locator3, alpha184_3_x_locator3);
  gfmult gfm_alpha185_0_x_locator0(10'b0000000001, locator0, alpha185_0_x_locator0);
  gfmult gfm_alpha185_1_x_locator1(10'b0101101011, locator1, alpha185_1_x_locator1);
  gfmult gfm_alpha185_2_x_locator2(10'b1000101000, locator2, alpha185_2_x_locator2);
  gfmult gfm_alpha185_3_x_locator3(10'b0101101101, locator3, alpha185_3_x_locator3);
  gfmult gfm_alpha186_0_x_locator0(10'b0000000001, locator0, alpha186_0_x_locator0);
  gfmult gfm_alpha186_1_x_locator1(10'b1010110001, locator1, alpha186_1_x_locator1);
  gfmult gfm_alpha186_2_x_locator2(10'b0010001010, locator2, alpha186_2_x_locator2);
  gfmult gfm_alpha186_3_x_locator3(10'b1010101000, locator3, alpha186_3_x_locator3);
  gfmult gfm_alpha187_0_x_locator0(10'b0000000001, locator0, alpha187_0_x_locator0);
  gfmult gfm_alpha187_1_x_locator1(10'b1101011100, locator1, alpha187_1_x_locator1);
  gfmult gfm_alpha187_2_x_locator2(10'b1000100110, locator2, alpha187_2_x_locator2);
  gfmult gfm_alpha187_3_x_locator3(10'b0001010101, locator3, alpha187_3_x_locator3);
  gfmult gfm_alpha188_0_x_locator0(10'b0000000001, locator0, alpha188_0_x_locator0);
  gfmult gfm_alpha188_1_x_locator1(10'b0110101110, locator1, alpha188_1_x_locator1);
  gfmult gfm_alpha188_2_x_locator2(10'b1010001101, locator2, alpha188_2_x_locator2);
  gfmult gfm_alpha188_3_x_locator3(10'b1010001111, locator3, alpha188_3_x_locator3);
  gfmult gfm_alpha189_0_x_locator0(10'b0000000001, locator0, alpha189_0_x_locator0);
  gfmult gfm_alpha189_1_x_locator1(10'b0011010111, locator1, alpha189_1_x_locator1);
  gfmult gfm_alpha189_2_x_locator2(10'b0110100001, locator2, alpha189_2_x_locator2);
  gfmult gfm_alpha189_3_x_locator3(10'b1111010110, locator3, alpha189_3_x_locator3);
  gfmult gfm_alpha190_0_x_locator0(10'b0000000001, locator0, alpha190_0_x_locator0);
  gfmult gfm_alpha190_1_x_locator1(10'b1001101111, locator1, alpha190_1_x_locator1);
  gfmult gfm_alpha190_2_x_locator2(10'b0101101010, locator2, alpha190_2_x_locator2);
  gfmult gfm_alpha190_3_x_locator3(10'b1101111100, locator3, alpha190_3_x_locator3);
  gfmult gfm_alpha191_0_x_locator0(10'b0000000001, locator0, alpha191_0_x_locator0);
  gfmult gfm_alpha191_1_x_locator1(10'b1100110011, locator1, alpha191_1_x_locator1);
  gfmult gfm_alpha191_2_x_locator2(10'b1001011110, locator2, alpha191_2_x_locator2);
  gfmult gfm_alpha191_3_x_locator3(10'b1001101011, locator3, alpha191_3_x_locator3);
  gfmult gfm_alpha192_0_x_locator0(10'b0000000001, locator0, alpha192_0_x_locator0);
  gfmult gfm_alpha192_1_x_locator1(10'b1110011101, locator1, alpha192_1_x_locator1);
  gfmult gfm_alpha192_2_x_locator2(10'b1010010011, locator2, alpha192_2_x_locator2);
  gfmult gfm_alpha192_3_x_locator3(10'b0111001110, locator3, alpha192_3_x_locator3);
  gfmult gfm_alpha193_0_x_locator0(10'b0000000001, locator0, alpha193_0_x_locator0);
  gfmult gfm_alpha193_1_x_locator1(10'b1111001010, locator1, alpha193_1_x_locator1);
  gfmult gfm_alpha193_2_x_locator2(10'b1110100010, locator2, alpha193_2_x_locator2);
  gfmult gfm_alpha193_3_x_locator3(10'b1100111111, locator3, alpha193_3_x_locator3);
  gfmult gfm_alpha194_0_x_locator0(10'b0000000001, locator0, alpha194_0_x_locator0);
  gfmult gfm_alpha194_1_x_locator1(10'b0111100101, locator1, alpha194_1_x_locator1);
  gfmult gfm_alpha194_2_x_locator2(10'b1011101100, locator2, alpha194_2_x_locator2);
  gfmult gfm_alpha194_3_x_locator3(10'b1111100000, locator3, alpha194_3_x_locator3);
  gfmult gfm_alpha195_0_x_locator0(10'b0000000001, locator0, alpha195_0_x_locator0);
  gfmult gfm_alpha195_1_x_locator1(10'b1011110110, locator1, alpha195_1_x_locator1);
  gfmult gfm_alpha195_2_x_locator2(10'b0010111011, locator2, alpha195_2_x_locator2);
  gfmult gfm_alpha195_3_x_locator3(10'b0001111100, locator3, alpha195_3_x_locator3);
  gfmult gfm_alpha196_0_x_locator0(10'b0000000001, locator0, alpha196_0_x_locator0);
  gfmult gfm_alpha196_1_x_locator1(10'b0101111011, locator1, alpha196_1_x_locator1);
  gfmult gfm_alpha196_2_x_locator2(10'b1100101000, locator2, alpha196_2_x_locator2);
  gfmult gfm_alpha196_3_x_locator3(10'b1000001011, locator3, alpha196_3_x_locator3);
  gfmult gfm_alpha197_0_x_locator0(10'b0000000001, locator0, alpha197_0_x_locator0);
  gfmult gfm_alpha197_1_x_locator1(10'b1010111001, locator1, alpha197_1_x_locator1);
  gfmult gfm_alpha197_2_x_locator2(10'b0011001010, locator2, alpha197_2_x_locator2);
  gfmult gfm_alpha197_3_x_locator3(10'b0111000010, locator3, alpha197_3_x_locator3);
  gfmult gfm_alpha198_0_x_locator0(10'b0000000001, locator0, alpha198_0_x_locator0);
  gfmult gfm_alpha198_1_x_locator1(10'b1101011000, locator1, alpha198_1_x_locator1);
  gfmult gfm_alpha198_2_x_locator2(10'b1000110110, locator2, alpha198_2_x_locator2);
  gfmult gfm_alpha198_3_x_locator3(10'b0100111010, locator3, alpha198_3_x_locator3);
  gfmult gfm_alpha199_0_x_locator0(10'b0000000001, locator0, alpha199_0_x_locator0);
  gfmult gfm_alpha199_1_x_locator1(10'b0110101100, locator1, alpha199_1_x_locator1);
  gfmult gfm_alpha199_2_x_locator2(10'b1010001001, locator2, alpha199_2_x_locator2);
  gfmult gfm_alpha199_3_x_locator3(10'b0100100101, locator3, alpha199_3_x_locator3);
  gfmult gfm_alpha200_0_x_locator0(10'b0000000001, locator0, alpha200_0_x_locator0);
  gfmult gfm_alpha200_1_x_locator1(10'b0011010110, locator1, alpha200_1_x_locator1);
  gfmult gfm_alpha200_2_x_locator2(10'b0110100000, locator2, alpha200_2_x_locator2);
  gfmult gfm_alpha200_3_x_locator3(10'b1010100001, locator3, alpha200_3_x_locator3);
  gfmult gfm_alpha201_0_x_locator0(10'b0000000001, locator0, alpha201_0_x_locator0);
  gfmult gfm_alpha201_1_x_locator1(10'b0001101011, locator1, alpha201_1_x_locator1);
  gfmult gfm_alpha201_2_x_locator2(10'b0001101000, locator2, alpha201_2_x_locator2);
  gfmult gfm_alpha201_3_x_locator3(10'b0011010101, locator3, alpha201_3_x_locator3);
  gfmult gfm_alpha202_0_x_locator0(10'b0000000001, locator0, alpha202_0_x_locator0);
  gfmult gfm_alpha202_1_x_locator1(10'b1000110001, locator1, alpha202_1_x_locator1);
  gfmult gfm_alpha202_2_x_locator2(10'b0000011010, locator2, alpha202_2_x_locator2);
  gfmult gfm_alpha202_3_x_locator3(10'b1010011111, locator3, alpha202_3_x_locator3);
  gfmult gfm_alpha203_0_x_locator0(10'b0000000001, locator0, alpha203_0_x_locator0);
  gfmult gfm_alpha203_1_x_locator1(10'b1100011100, locator1, alpha203_1_x_locator1);
  gfmult gfm_alpha203_2_x_locator2(10'b1000000010, locator2, alpha203_2_x_locator2);
  gfmult gfm_alpha203_3_x_locator3(10'b1111010100, locator3, alpha203_3_x_locator3);
  gfmult gfm_alpha204_0_x_locator0(10'b0000000001, locator0, alpha204_0_x_locator0);
  gfmult gfm_alpha204_1_x_locator1(10'b0110001110, locator1, alpha204_1_x_locator1);
  gfmult gfm_alpha204_2_x_locator2(10'b1010000100, locator2, alpha204_2_x_locator2);
  gfmult gfm_alpha204_3_x_locator3(10'b1001111110, locator3, alpha204_3_x_locator3);
  gfmult gfm_alpha205_0_x_locator0(10'b0000000001, locator0, alpha205_0_x_locator0);
  gfmult gfm_alpha205_1_x_locator1(10'b0011000111, locator1, alpha205_1_x_locator1);
  gfmult gfm_alpha205_2_x_locator2(10'b0010100001, locator2, alpha205_2_x_locator2);
  gfmult gfm_alpha205_3_x_locator3(10'b1101001001, locator3, alpha205_3_x_locator3);
  gfmult gfm_alpha206_0_x_locator0(10'b0000000001, locator0, alpha206_0_x_locator0);
  gfmult gfm_alpha206_1_x_locator1(10'b1001100111, locator1, alpha206_1_x_locator1);
  gfmult gfm_alpha206_2_x_locator2(10'b0100101010, locator2, alpha206_2_x_locator2);
  gfmult gfm_alpha206_3_x_locator3(10'b0011101000, locator3, alpha206_3_x_locator3);
  gfmult gfm_alpha207_0_x_locator0(10'b0000000001, locator0, alpha207_0_x_locator0);
  gfmult gfm_alpha207_1_x_locator1(10'b1100110111, locator1, alpha207_1_x_locator1);
  gfmult gfm_alpha207_2_x_locator2(10'b1001001110, locator2, alpha207_2_x_locator2);
  gfmult gfm_alpha207_3_x_locator3(10'b0000011101, locator3, alpha207_3_x_locator3);
  gfmult gfm_alpha208_0_x_locator0(10'b0000000001, locator0, alpha208_0_x_locator0);
  gfmult gfm_alpha208_1_x_locator1(10'b1110011111, locator1, alpha208_1_x_locator1);
  gfmult gfm_alpha208_2_x_locator2(10'b1010010111, locator2, alpha208_2_x_locator2);
  gfmult gfm_alpha208_3_x_locator3(10'b1010000110, locator3, alpha208_3_x_locator3);
  gfmult gfm_alpha209_0_x_locator0(10'b0000000001, locator0, alpha209_0_x_locator0);
  gfmult gfm_alpha209_1_x_locator1(10'b1111001011, locator1, alpha209_1_x_locator1);
  gfmult gfm_alpha209_2_x_locator2(10'b1110100011, locator2, alpha209_2_x_locator2);
  gfmult gfm_alpha209_3_x_locator3(10'b1101010110, locator3, alpha209_3_x_locator3);
  gfmult gfm_alpha210_0_x_locator0(10'b0000000001, locator0, alpha210_0_x_locator0);
  gfmult gfm_alpha210_1_x_locator1(10'b1111100001, locator1, alpha210_1_x_locator1);
  gfmult gfm_alpha210_2_x_locator2(10'b1111101110, locator2, alpha210_2_x_locator2);
  gfmult gfm_alpha210_3_x_locator3(10'b1101101100, locator3, alpha210_3_x_locator3);
  gfmult gfm_alpha211_0_x_locator0(10'b0000000001, locator0, alpha211_0_x_locator0);
  gfmult gfm_alpha211_1_x_locator1(10'b1111110100, locator1, alpha211_1_x_locator1);
  gfmult gfm_alpha211_2_x_locator2(10'b1011111111, locator2, alpha211_2_x_locator2);
  gfmult gfm_alpha211_3_x_locator3(10'b1001101001, locator3, alpha211_3_x_locator3);
  gfmult gfm_alpha212_0_x_locator0(10'b0000000001, locator0, alpha212_0_x_locator0);
  gfmult gfm_alpha212_1_x_locator1(10'b0111111010, locator1, alpha212_1_x_locator1);
  gfmult gfm_alpha212_2_x_locator2(10'b1110111001, locator2, alpha212_2_x_locator2);
  gfmult gfm_alpha212_3_x_locator3(10'b0011001100, locator3, alpha212_3_x_locator3);
  gfmult gfm_alpha213_0_x_locator0(10'b0000000001, locator0, alpha213_0_x_locator0);
  gfmult gfm_alpha213_1_x_locator1(10'b0011111101, locator1, alpha213_1_x_locator1);
  gfmult gfm_alpha213_2_x_locator2(10'b0111101100, locator2, alpha213_2_x_locator2);
  gfmult gfm_alpha213_3_x_locator3(10'b1000011101, locator3, alpha213_3_x_locator3);
  gfmult gfm_alpha214_0_x_locator0(10'b0000000001, locator0, alpha214_0_x_locator0);
  gfmult gfm_alpha214_1_x_locator1(10'b1001111010, locator1, alpha214_1_x_locator1);
  gfmult gfm_alpha214_2_x_locator2(10'b0001111011, locator2, alpha214_2_x_locator2);
  gfmult gfm_alpha214_3_x_locator3(10'b1011000110, locator3, alpha214_3_x_locator3);
  gfmult gfm_alpha215_0_x_locator0(10'b0000000001, locator0, alpha215_0_x_locator0);
  gfmult gfm_alpha215_1_x_locator1(10'b0100111101, locator1, alpha215_1_x_locator1);
  gfmult gfm_alpha215_2_x_locator2(10'b1100011000, locator2, alpha215_2_x_locator2);
  gfmult gfm_alpha215_3_x_locator3(10'b1101011110, locator3, alpha215_3_x_locator3);
  gfmult gfm_alpha216_0_x_locator0(10'b0000000001, locator0, alpha216_0_x_locator0);
  gfmult gfm_alpha216_1_x_locator1(10'b1010011010, locator1, alpha216_1_x_locator1);
  gfmult gfm_alpha216_2_x_locator2(10'b0011000110, locator2, alpha216_2_x_locator2);
  gfmult gfm_alpha216_3_x_locator3(10'b1101101101, locator3, alpha216_3_x_locator3);
  gfmult gfm_alpha217_0_x_locator0(10'b0000000001, locator0, alpha217_0_x_locator0);
  gfmult gfm_alpha217_1_x_locator1(10'b0101001101, locator1, alpha217_1_x_locator1);
  gfmult gfm_alpha217_2_x_locator2(10'b1000110101, locator2, alpha217_2_x_locator2);
  gfmult gfm_alpha217_3_x_locator3(10'b1011101000, locator3, alpha217_3_x_locator3);
  gfmult gfm_alpha218_0_x_locator0(10'b0000000001, locator0, alpha218_0_x_locator0);
  gfmult gfm_alpha218_1_x_locator1(10'b1010100010, locator1, alpha218_1_x_locator1);
  gfmult gfm_alpha218_2_x_locator2(10'b0110001111, locator2, alpha218_2_x_locator2);
  gfmult gfm_alpha218_3_x_locator3(10'b0001011101, locator3, alpha218_3_x_locator3);
  gfmult gfm_alpha219_0_x_locator0(10'b0000000001, locator0, alpha219_0_x_locator0);
  gfmult gfm_alpha219_1_x_locator1(10'b0101010001, locator1, alpha219_1_x_locator1);
  gfmult gfm_alpha219_2_x_locator2(10'b1101100101, locator2, alpha219_2_x_locator2);
  gfmult gfm_alpha219_3_x_locator3(10'b1010001110, locator3, alpha219_3_x_locator3);
  gfmult gfm_alpha220_0_x_locator0(10'b0000000001, locator0, alpha220_0_x_locator0);
  gfmult gfm_alpha220_1_x_locator1(10'b1010101100, locator1, alpha220_1_x_locator1);
  gfmult gfm_alpha220_2_x_locator2(10'b0111011011, locator2, alpha220_2_x_locator2);
  gfmult gfm_alpha220_3_x_locator3(10'b1101010111, locator3, alpha220_3_x_locator3);
  gfmult gfm_alpha221_0_x_locator0(10'b0000000001, locator0, alpha221_0_x_locator0);
  gfmult gfm_alpha221_1_x_locator1(10'b0101010110, locator1, alpha221_1_x_locator1);
  gfmult gfm_alpha221_2_x_locator2(10'b1101110000, locator2, alpha221_2_x_locator2);
  gfmult gfm_alpha221_3_x_locator3(10'b1111101101, locator3, alpha221_3_x_locator3);
  gfmult gfm_alpha222_0_x_locator0(10'b0000000001, locator0, alpha222_0_x_locator0);
  gfmult gfm_alpha222_1_x_locator1(10'b0010101011, locator1, alpha222_1_x_locator1);
  gfmult gfm_alpha222_2_x_locator2(10'b0011011100, locator2, alpha222_2_x_locator2);
  gfmult gfm_alpha222_3_x_locator3(10'b1011111000, locator3, alpha222_3_x_locator3);
  gfmult gfm_alpha223_0_x_locator0(10'b0000000001, locator0, alpha223_0_x_locator0);
  gfmult gfm_alpha223_1_x_locator1(10'b1001010001, locator1, alpha223_1_x_locator1);
  gfmult gfm_alpha223_2_x_locator2(10'b0000110111, locator2, alpha223_2_x_locator2);
  gfmult gfm_alpha223_3_x_locator3(10'b0001011111, locator3, alpha223_3_x_locator3);
  gfmult gfm_alpha224_0_x_locator0(10'b0000000001, locator0, alpha224_0_x_locator0);
  gfmult gfm_alpha224_1_x_locator1(10'b1100101100, locator1, alpha224_1_x_locator1);
  gfmult gfm_alpha224_2_x_locator2(10'b1100001011, locator2, alpha224_2_x_locator2);
  gfmult gfm_alpha224_3_x_locator3(10'b1110001100, locator3, alpha224_3_x_locator3);
  gfmult gfm_alpha225_0_x_locator0(10'b0000000001, locator0, alpha225_0_x_locator0);
  gfmult gfm_alpha225_1_x_locator1(10'b0110010110, locator1, alpha225_1_x_locator1);
  gfmult gfm_alpha225_2_x_locator2(10'b1111000100, locator2, alpha225_2_x_locator2);
  gfmult gfm_alpha225_3_x_locator3(10'b1001110101, locator3, alpha225_3_x_locator3);
  gfmult gfm_alpha226_0_x_locator0(10'b0000000001, locator0, alpha226_0_x_locator0);
  gfmult gfm_alpha226_1_x_locator1(10'b0011001011, locator1, alpha226_1_x_locator1);
  gfmult gfm_alpha226_2_x_locator2(10'b0011110001, locator2, alpha226_2_x_locator2);
  gfmult gfm_alpha226_3_x_locator3(10'b1011001011, locator3, alpha226_3_x_locator3);
  gfmult gfm_alpha227_0_x_locator0(10'b0000000001, locator0, alpha227_0_x_locator0);
  gfmult gfm_alpha227_1_x_locator1(10'b1001100001, locator1, alpha227_1_x_locator1);
  gfmult gfm_alpha227_2_x_locator2(10'b0100111110, locator2, alpha227_2_x_locator2);
  gfmult gfm_alpha227_3_x_locator3(10'b0111011010, locator3, alpha227_3_x_locator3);
  gfmult gfm_alpha228_0_x_locator0(10'b0000000001, locator0, alpha228_0_x_locator0);
  gfmult gfm_alpha228_1_x_locator1(10'b1100110100, locator1, alpha228_1_x_locator1);
  gfmult gfm_alpha228_2_x_locator2(10'b1001001011, locator2, alpha228_2_x_locator2);
  gfmult gfm_alpha228_3_x_locator3(10'b0100111001, locator3, alpha228_3_x_locator3);
  gfmult gfm_alpha229_0_x_locator0(10'b0000000001, locator0, alpha229_0_x_locator0);
  gfmult gfm_alpha229_1_x_locator1(10'b0110011010, locator1, alpha229_1_x_locator1);
  gfmult gfm_alpha229_2_x_locator2(10'b1110010100, locator2, alpha229_2_x_locator2);
  gfmult gfm_alpha229_3_x_locator3(10'b0010100110, locator3, alpha229_3_x_locator3);
  gfmult gfm_alpha230_0_x_locator0(10'b0000000001, locator0, alpha230_0_x_locator0);
  gfmult gfm_alpha230_1_x_locator1(10'b0011001101, locator1, alpha230_1_x_locator1);
  gfmult gfm_alpha230_2_x_locator2(10'b0011100101, locator2, alpha230_2_x_locator2);
  gfmult gfm_alpha230_3_x_locator3(10'b1100010010, locator3, alpha230_3_x_locator3);
  gfmult gfm_alpha231_0_x_locator0(10'b0000000001, locator0, alpha231_0_x_locator0);
  gfmult gfm_alpha231_1_x_locator1(10'b1001100010, locator1, alpha231_1_x_locator1);
  gfmult gfm_alpha231_2_x_locator2(10'b0100111011, locator2, alpha231_2_x_locator2);
  gfmult gfm_alpha231_3_x_locator3(10'b0101100000, locator3, alpha231_3_x_locator3);
  gfmult gfm_alpha232_0_x_locator0(10'b0000000001, locator0, alpha232_0_x_locator0);
  gfmult gfm_alpha232_1_x_locator1(10'b0100110001, locator1, alpha232_1_x_locator1);
  gfmult gfm_alpha232_2_x_locator2(10'b1101001000, locator2, alpha232_2_x_locator2);
  gfmult gfm_alpha232_3_x_locator3(10'b0000101100, locator3, alpha232_3_x_locator3);
  gfmult gfm_alpha233_0_x_locator0(10'b0000000001, locator0, alpha233_0_x_locator0);
  gfmult gfm_alpha233_1_x_locator1(10'b1010011100, locator1, alpha233_1_x_locator1);
  gfmult gfm_alpha233_2_x_locator2(10'b0011010010, locator2, alpha233_2_x_locator2);
  gfmult gfm_alpha233_3_x_locator3(10'b1000000001, locator3, alpha233_3_x_locator3);
  gfmult gfm_alpha234_0_x_locator0(10'b0000000001, locator0, alpha234_0_x_locator0);
  gfmult gfm_alpha234_1_x_locator1(10'b0101001110, locator1, alpha234_1_x_locator1);
  gfmult gfm_alpha234_2_x_locator2(10'b1000110000, locator2, alpha234_2_x_locator2);
  gfmult gfm_alpha234_3_x_locator3(10'b0011000001, locator3, alpha234_3_x_locator3);
  gfmult gfm_alpha235_0_x_locator0(10'b0000000001, locator0, alpha235_0_x_locator0);
  gfmult gfm_alpha235_1_x_locator1(10'b0010100111, locator1, alpha235_1_x_locator1);
  gfmult gfm_alpha235_2_x_locator2(10'b0010001100, locator2, alpha235_2_x_locator2);
  gfmult gfm_alpha235_3_x_locator3(10'b0010011001, locator3, alpha235_3_x_locator3);
  gfmult gfm_alpha236_0_x_locator0(10'b0000000001, locator0, alpha236_0_x_locator0);
  gfmult gfm_alpha236_1_x_locator1(10'b1001010111, locator1, alpha236_1_x_locator1);
  gfmult gfm_alpha236_2_x_locator2(10'b0000100011, locator2, alpha236_2_x_locator2);
  gfmult gfm_alpha236_3_x_locator3(10'b0010010010, locator3, alpha236_3_x_locator3);
  gfmult gfm_alpha237_0_x_locator0(10'b0000000001, locator0, alpha237_0_x_locator0);
  gfmult gfm_alpha237_1_x_locator1(10'b1100101111, locator1, alpha237_1_x_locator1);
  gfmult gfm_alpha237_2_x_locator2(10'b1100001110, locator2, alpha237_2_x_locator2);
  gfmult gfm_alpha237_3_x_locator3(10'b0100010000, locator3, alpha237_3_x_locator3);
  gfmult gfm_alpha238_0_x_locator0(10'b0000000001, locator0, alpha238_0_x_locator0);
  gfmult gfm_alpha238_1_x_locator1(10'b1110010011, locator1, alpha238_1_x_locator1);
  gfmult gfm_alpha238_2_x_locator2(10'b1011000111, locator2, alpha238_2_x_locator2);
  gfmult gfm_alpha238_3_x_locator3(10'b0000100010, locator3, alpha238_3_x_locator3);
  gfmult gfm_alpha239_0_x_locator0(10'b0000000001, locator0, alpha239_0_x_locator0);
  gfmult gfm_alpha239_1_x_locator1(10'b1111001101, locator1, alpha239_1_x_locator1);
  gfmult gfm_alpha239_2_x_locator2(10'b1110110111, locator2, alpha239_2_x_locator2);
  gfmult gfm_alpha239_3_x_locator3(10'b0100000110, locator3, alpha239_3_x_locator3);
  gfmult gfm_alpha240_0_x_locator0(10'b0000000001, locator0, alpha240_0_x_locator0);
  gfmult gfm_alpha240_1_x_locator1(10'b1111100010, locator1, alpha240_1_x_locator1);
  gfmult gfm_alpha240_2_x_locator2(10'b1111101011, locator2, alpha240_2_x_locator2);
  gfmult gfm_alpha240_3_x_locator3(10'b1100100110, locator3, alpha240_3_x_locator3);
  gfmult gfm_alpha241_0_x_locator0(10'b0000000001, locator0, alpha241_0_x_locator0);
  gfmult gfm_alpha241_1_x_locator1(10'b0111110001, locator1, alpha241_1_x_locator1);
  gfmult gfm_alpha241_2_x_locator2(10'b1111111100, locator2, alpha241_2_x_locator2);
  gfmult gfm_alpha241_3_x_locator3(10'b1101100010, locator3, alpha241_3_x_locator3);
  gfmult gfm_alpha242_0_x_locator0(10'b0000000001, locator0, alpha242_0_x_locator0);
  gfmult gfm_alpha242_1_x_locator1(10'b1011111100, locator1, alpha242_1_x_locator1);
  gfmult gfm_alpha242_2_x_locator2(10'b0011111111, locator2, alpha242_2_x_locator2);
  gfmult gfm_alpha242_3_x_locator3(10'b0101101110, locator3, alpha242_3_x_locator3);
  gfmult gfm_alpha243_0_x_locator0(10'b0000000001, locator0, alpha243_0_x_locator0);
  gfmult gfm_alpha243_1_x_locator1(10'b0101111110, locator1, alpha243_1_x_locator1);
  gfmult gfm_alpha243_2_x_locator2(10'b1100111001, locator2, alpha243_2_x_locator2);
  gfmult gfm_alpha243_3_x_locator3(10'b1100101011, locator3, alpha243_3_x_locator3);
  gfmult gfm_alpha244_0_x_locator0(10'b0000000001, locator0, alpha244_0_x_locator0);
  gfmult gfm_alpha244_1_x_locator1(10'b0010111111, locator1, alpha244_1_x_locator1);
  gfmult gfm_alpha244_2_x_locator2(10'b0111001100, locator2, alpha244_2_x_locator2);
  gfmult gfm_alpha244_3_x_locator3(10'b0111100110, locator3, alpha244_3_x_locator3);
  gfmult gfm_alpha245_0_x_locator0(10'b0000000001, locator0, alpha245_0_x_locator0);
  gfmult gfm_alpha245_1_x_locator1(10'b1001011011, locator1, alpha245_1_x_locator1);
  gfmult gfm_alpha245_2_x_locator2(10'b0001110011, locator2, alpha245_2_x_locator2);
  gfmult gfm_alpha245_3_x_locator3(10'b1100111010, locator3, alpha245_3_x_locator3);
  gfmult gfm_alpha246_0_x_locator0(10'b0000000001, locator0, alpha246_0_x_locator0);
  gfmult gfm_alpha246_1_x_locator1(10'b1100101001, locator1, alpha246_1_x_locator1);
  gfmult gfm_alpha246_2_x_locator2(10'b1100011010, locator2, alpha246_2_x_locator2);
  gfmult gfm_alpha246_3_x_locator3(10'b0101100101, locator3, alpha246_3_x_locator3);
  gfmult gfm_alpha247_0_x_locator0(10'b0000000001, locator0, alpha247_0_x_locator0);
  gfmult gfm_alpha247_1_x_locator1(10'b1110010000, locator1, alpha247_1_x_locator1);
  gfmult gfm_alpha247_2_x_locator2(10'b1011000010, locator2, alpha247_2_x_locator2);
  gfmult gfm_alpha247_3_x_locator3(10'b1010101001, locator3, alpha247_3_x_locator3);
  gfmult gfm_alpha248_0_x_locator0(10'b0000000001, locator0, alpha248_0_x_locator0);
  gfmult gfm_alpha248_1_x_locator1(10'b0111001000, locator1, alpha248_1_x_locator1);
  gfmult gfm_alpha248_2_x_locator2(10'b1010110100, locator2, alpha248_2_x_locator2);
  gfmult gfm_alpha248_3_x_locator3(10'b0011010100, locator3, alpha248_3_x_locator3);
  gfmult gfm_alpha249_0_x_locator0(10'b0000000001, locator0, alpha249_0_x_locator0);
  gfmult gfm_alpha249_1_x_locator1(10'b0011100100, locator1, alpha249_1_x_locator1);
  gfmult gfm_alpha249_2_x_locator2(10'b0010101101, locator2, alpha249_2_x_locator2);
  gfmult gfm_alpha249_3_x_locator3(10'b1000011110, locator3, alpha249_3_x_locator3);
  gfmult gfm_alpha250_0_x_locator0(10'b0000000001, locator0, alpha250_0_x_locator0);
  gfmult gfm_alpha250_1_x_locator1(10'b0001110010, locator1, alpha250_1_x_locator1);
  gfmult gfm_alpha250_2_x_locator2(10'b0100101001, locator2, alpha250_2_x_locator2);
  gfmult gfm_alpha250_3_x_locator3(10'b1101000101, locator3, alpha250_3_x_locator3);
  gfmult gfm_alpha251_0_x_locator0(10'b0000000001, locator0, alpha251_0_x_locator0);
  gfmult gfm_alpha251_1_x_locator1(10'b0000111001, locator1, alpha251_1_x_locator1);
  gfmult gfm_alpha251_2_x_locator2(10'b0101001000, locator2, alpha251_2_x_locator2);
  gfmult gfm_alpha251_3_x_locator3(10'b1011101101, locator3, alpha251_3_x_locator3);
  gfmult gfm_alpha252_0_x_locator0(10'b0000000001, locator0, alpha252_0_x_locator0);
  gfmult gfm_alpha252_1_x_locator1(10'b1000011000, locator1, alpha252_1_x_locator1);
  gfmult gfm_alpha252_2_x_locator2(10'b0001010010, locator2, alpha252_2_x_locator2);
  gfmult gfm_alpha252_3_x_locator3(10'b1011011000, locator3, alpha252_3_x_locator3);
  gfmult gfm_alpha253_0_x_locator0(10'b0000000001, locator0, alpha253_0_x_locator0);
  gfmult gfm_alpha253_1_x_locator1(10'b0100001100, locator1, alpha253_1_x_locator1);
  gfmult gfm_alpha253_2_x_locator2(10'b1000010000, locator2, alpha253_2_x_locator2);
  gfmult gfm_alpha253_3_x_locator3(10'b0001011011, locator3, alpha253_3_x_locator3);
  gfmult gfm_alpha254_0_x_locator0(10'b0000000001, locator0, alpha254_0_x_locator0);
  gfmult gfm_alpha254_1_x_locator1(10'b0010000110, locator1, alpha254_1_x_locator1);
  gfmult gfm_alpha254_2_x_locator2(10'b0010000100, locator2, alpha254_2_x_locator2);
  gfmult gfm_alpha254_3_x_locator3(10'b0110001000, locator3, alpha254_3_x_locator3);
  gfmult gfm_alpha255_0_x_locator0(10'b0000000001, locator0, alpha255_0_x_locator0);
  gfmult gfm_alpha255_1_x_locator1(10'b0001000011, locator1, alpha255_1_x_locator1);
  gfmult gfm_alpha255_2_x_locator2(10'b0000100001, locator2, alpha255_2_x_locator2);
  gfmult gfm_alpha255_3_x_locator3(10'b0000110001, locator3, alpha255_3_x_locator3);
  gfmult gfm_alpha256_0_x_locator0(10'b0000000001, locator0, alpha256_0_x_locator0);
  gfmult gfm_alpha256_1_x_locator1(10'b1000100101, locator1, alpha256_1_x_locator1);
  gfmult gfm_alpha256_2_x_locator2(10'b0100001010, locator2, alpha256_2_x_locator2);
  gfmult gfm_alpha256_3_x_locator3(10'b0010000111, locator3, alpha256_3_x_locator3);
  gfmult gfm_alpha257_0_x_locator0(10'b0000000001, locator0, alpha257_0_x_locator0);
  gfmult gfm_alpha257_1_x_locator1(10'b1100010110, locator1, alpha257_1_x_locator1);
  gfmult gfm_alpha257_2_x_locator2(10'b1001000110, locator2, alpha257_2_x_locator2);
  gfmult gfm_alpha257_3_x_locator3(10'b1110010111, locator3, alpha257_3_x_locator3);
  gfmult gfm_alpha258_0_x_locator0(10'b0000000001, locator0, alpha258_0_x_locator0);
  gfmult gfm_alpha258_1_x_locator1(10'b0110001011, locator1, alpha258_1_x_locator1);
  gfmult gfm_alpha258_2_x_locator2(10'b1010010101, locator2, alpha258_2_x_locator2);
  gfmult gfm_alpha258_3_x_locator3(10'b1111110101, locator3, alpha258_3_x_locator3);
  gfmult gfm_alpha259_0_x_locator0(10'b0000000001, locator0, alpha259_0_x_locator0);
  gfmult gfm_alpha259_1_x_locator1(10'b1011000001, locator1, alpha259_1_x_locator1);
  gfmult gfm_alpha259_2_x_locator2(10'b0110100111, locator2, alpha259_2_x_locator2);
  gfmult gfm_alpha259_3_x_locator3(10'b1011111011, locator3, alpha259_3_x_locator3);
  gfmult gfm_alpha260_0_x_locator0(10'b0000000001, locator0, alpha260_0_x_locator0);
  gfmult gfm_alpha260_1_x_locator1(10'b1101100100, locator1, alpha260_1_x_locator1);
  gfmult gfm_alpha260_2_x_locator2(10'b1101101111, locator2, alpha260_2_x_locator2);
  gfmult gfm_alpha260_3_x_locator3(10'b0111011100, locator3, alpha260_3_x_locator3);
  gfmult gfm_alpha261_0_x_locator0(10'b0000000001, locator0, alpha261_0_x_locator0);
  gfmult gfm_alpha261_1_x_locator1(10'b0110110010, locator1, alpha261_1_x_locator1);
  gfmult gfm_alpha261_2_x_locator2(10'b1111011101, locator2, alpha261_2_x_locator2);
  gfmult gfm_alpha261_3_x_locator3(10'b1000111111, locator3, alpha261_3_x_locator3);
  gfmult gfm_alpha262_0_x_locator0(10'b0000000001, locator0, alpha262_0_x_locator0);
  gfmult gfm_alpha262_1_x_locator1(10'b0011011001, locator1, alpha262_1_x_locator1);
  gfmult gfm_alpha262_2_x_locator2(10'b0111110101, locator2, alpha262_2_x_locator2);
  gfmult gfm_alpha262_3_x_locator3(10'b1111000000, locator3, alpha262_3_x_locator3);
  gfmult gfm_alpha263_0_x_locator0(10'b0000000001, locator0, alpha263_0_x_locator0);
  gfmult gfm_alpha263_1_x_locator1(10'b1001101000, locator1, alpha263_1_x_locator1);
  gfmult gfm_alpha263_2_x_locator2(10'b0101111111, locator2, alpha263_2_x_locator2);
  gfmult gfm_alpha263_3_x_locator3(10'b0001111000, locator3, alpha263_3_x_locator3);
  gfmult gfm_alpha264_0_x_locator0(10'b0000000001, locator0, alpha264_0_x_locator0);
  gfmult gfm_alpha264_1_x_locator1(10'b0100110100, locator1, alpha264_1_x_locator1);
  gfmult gfm_alpha264_2_x_locator2(10'b1101011001, locator2, alpha264_2_x_locator2);
  gfmult gfm_alpha264_3_x_locator3(10'b0000001111, locator3, alpha264_3_x_locator3);
  gfmult gfm_alpha265_0_x_locator0(10'b0000000001, locator0, alpha265_0_x_locator0);
  gfmult gfm_alpha265_1_x_locator1(10'b0010011010, locator1, alpha265_1_x_locator1);
  gfmult gfm_alpha265_2_x_locator2(10'b0111010100, locator2, alpha265_2_x_locator2);
  gfmult gfm_alpha265_3_x_locator3(10'b1110000110, locator3, alpha265_3_x_locator3);
  gfmult gfm_alpha266_0_x_locator0(10'b0000000001, locator0, alpha266_0_x_locator0);
  gfmult gfm_alpha266_1_x_locator1(10'b0001001101, locator1, alpha266_1_x_locator1);
  gfmult gfm_alpha266_2_x_locator2(10'b0001110101, locator2, alpha266_2_x_locator2);
  gfmult gfm_alpha266_3_x_locator3(10'b1101110110, locator3, alpha266_3_x_locator3);
  gfmult gfm_alpha267_0_x_locator0(10'b0000000001, locator0, alpha267_0_x_locator0);
  gfmult gfm_alpha267_1_x_locator1(10'b1000100010, locator1, alpha267_1_x_locator1);
  gfmult gfm_alpha267_2_x_locator2(10'b0100011111, locator2, alpha267_2_x_locator2);
  gfmult gfm_alpha267_3_x_locator3(10'b1101101000, locator3, alpha267_3_x_locator3);
  gfmult gfm_alpha268_0_x_locator0(10'b0000000001, locator0, alpha268_0_x_locator0);
  gfmult gfm_alpha268_1_x_locator1(10'b0100010001, locator1, alpha268_1_x_locator1);
  gfmult gfm_alpha268_2_x_locator2(10'b1101000001, locator2, alpha268_2_x_locator2);
  gfmult gfm_alpha268_3_x_locator3(10'b0001101101, locator3, alpha268_3_x_locator3);
  gfmult gfm_alpha269_0_x_locator0(10'b0000000001, locator0, alpha269_0_x_locator0);
  gfmult gfm_alpha269_1_x_locator1(10'b1010001100, locator1, alpha269_1_x_locator1);
  gfmult gfm_alpha269_2_x_locator2(10'b0111010010, locator2, alpha269_2_x_locator2);
  gfmult gfm_alpha269_3_x_locator3(10'b1010001000, locator3, alpha269_3_x_locator3);
  gfmult gfm_alpha270_0_x_locator0(10'b0000000001, locator0, alpha270_0_x_locator0);
  gfmult gfm_alpha270_1_x_locator1(10'b0101000110, locator1, alpha270_1_x_locator1);
  gfmult gfm_alpha270_2_x_locator2(10'b1001110000, locator2, alpha270_2_x_locator2);
  gfmult gfm_alpha270_3_x_locator3(10'b0001010001, locator3, alpha270_3_x_locator3);
  gfmult gfm_alpha271_0_x_locator0(10'b0000000001, locator0, alpha271_0_x_locator0);
  gfmult gfm_alpha271_1_x_locator1(10'b0010100011, locator1, alpha271_1_x_locator1);
  gfmult gfm_alpha271_2_x_locator2(10'b0010011100, locator2, alpha271_2_x_locator2);
  gfmult gfm_alpha271_3_x_locator3(10'b0010001011, locator3, alpha271_3_x_locator3);
  gfmult gfm_alpha272_0_x_locator0(10'b0000000001, locator0, alpha272_0_x_locator0);
  gfmult gfm_alpha272_1_x_locator1(10'b1001010101, locator1, alpha272_1_x_locator1);
  gfmult gfm_alpha272_2_x_locator2(10'b0000100111, locator2, alpha272_2_x_locator2);
  gfmult gfm_alpha272_3_x_locator3(10'b0110010010, locator3, alpha272_3_x_locator3);
  gfmult gfm_alpha273_0_x_locator0(10'b0000000001, locator0, alpha273_0_x_locator0);
  gfmult gfm_alpha273_1_x_locator1(10'b1100101110, locator1, alpha273_1_x_locator1);
  gfmult gfm_alpha273_2_x_locator2(10'b1100001111, locator2, alpha273_2_x_locator2);
  gfmult gfm_alpha273_3_x_locator3(10'b0100110000, locator3, alpha273_3_x_locator3);
  gfmult gfm_alpha274_0_x_locator0(10'b0000000001, locator0, alpha274_0_x_locator0);
  gfmult gfm_alpha274_1_x_locator1(10'b0110010111, locator1, alpha274_1_x_locator1);
  gfmult gfm_alpha274_2_x_locator2(10'b1111000101, locator2, alpha274_2_x_locator2);
  gfmult gfm_alpha274_3_x_locator3(10'b0000100110, locator3, alpha274_3_x_locator3);
  gfmult gfm_alpha275_0_x_locator0(10'b0000000001, locator0, alpha275_0_x_locator0);
  gfmult gfm_alpha275_1_x_locator1(10'b1011001111, locator1, alpha275_1_x_locator1);
  gfmult gfm_alpha275_2_x_locator2(10'b0111110011, locator2, alpha275_2_x_locator2);
  gfmult gfm_alpha275_3_x_locator3(10'b1100000010, locator3, alpha275_3_x_locator3);
  gfmult gfm_alpha276_0_x_locator0(10'b0000000001, locator0, alpha276_0_x_locator0);
  gfmult gfm_alpha276_1_x_locator1(10'b1101100011, locator1, alpha276_1_x_locator1);
  gfmult gfm_alpha276_2_x_locator2(10'b1101111010, locator2, alpha276_2_x_locator2);
  gfmult gfm_alpha276_3_x_locator3(10'b0101100010, locator3, alpha276_3_x_locator3);
  gfmult gfm_alpha277_0_x_locator0(10'b0000000001, locator0, alpha277_0_x_locator0);
  gfmult gfm_alpha277_1_x_locator1(10'b1110110101, locator1, alpha277_1_x_locator1);
  gfmult gfm_alpha277_2_x_locator2(10'b1011011010, locator2, alpha277_2_x_locator2);
  gfmult gfm_alpha277_3_x_locator3(10'b0100101110, locator3, alpha277_3_x_locator3);
  gfmult gfm_alpha278_0_x_locator0(10'b0000000001, locator0, alpha278_0_x_locator0);
  gfmult gfm_alpha278_1_x_locator1(10'b1111011110, locator1, alpha278_1_x_locator1);
  gfmult gfm_alpha278_2_x_locator2(10'b1010110010, locator2, alpha278_2_x_locator2);
  gfmult gfm_alpha278_3_x_locator3(10'b1100100011, locator3, alpha278_3_x_locator3);
  gfmult gfm_alpha279_0_x_locator0(10'b0000000001, locator0, alpha279_0_x_locator0);
  gfmult gfm_alpha279_1_x_locator1(10'b0111101111, locator1, alpha279_1_x_locator1);
  gfmult gfm_alpha279_2_x_locator2(10'b1010101000, locator2, alpha279_2_x_locator2);
  gfmult gfm_alpha279_3_x_locator3(10'b0111100111, locator3, alpha279_3_x_locator3);
  gfmult gfm_alpha280_0_x_locator0(10'b0000000001, locator0, alpha280_0_x_locator0);
  gfmult gfm_alpha280_1_x_locator1(10'b1011110011, locator1, alpha280_1_x_locator1);
  gfmult gfm_alpha280_2_x_locator2(10'b0010101010, locator2, alpha280_2_x_locator2);
  gfmult gfm_alpha280_3_x_locator3(10'b1110111011, locator3, alpha280_3_x_locator3);
  gfmult gfm_alpha281_0_x_locator0(10'b0000000001, locator0, alpha281_0_x_locator0);
  gfmult gfm_alpha281_1_x_locator1(10'b1101111101, locator1, alpha281_1_x_locator1);
  gfmult gfm_alpha281_2_x_locator2(10'b1000101110, locator2, alpha281_2_x_locator2);
  gfmult gfm_alpha281_3_x_locator3(10'b0111110100, locator3, alpha281_3_x_locator3);
  gfmult gfm_alpha282_0_x_locator0(10'b0000000001, locator0, alpha282_0_x_locator0);
  gfmult gfm_alpha282_1_x_locator1(10'b1110111010, locator1, alpha282_1_x_locator1);
  gfmult gfm_alpha282_2_x_locator2(10'b1010001111, locator2, alpha282_2_x_locator2);
  gfmult gfm_alpha282_3_x_locator3(10'b1000111010, locator3, alpha282_3_x_locator3);
  gfmult gfm_alpha283_0_x_locator0(10'b0000000001, locator0, alpha283_0_x_locator0);
  gfmult gfm_alpha283_1_x_locator1(10'b0111011101, locator1, alpha283_1_x_locator1);
  gfmult gfm_alpha283_2_x_locator2(10'b1110100101, locator2, alpha283_2_x_locator2);
  gfmult gfm_alpha283_3_x_locator3(10'b0101000101, locator3, alpha283_3_x_locator3);
  gfmult gfm_alpha284_0_x_locator0(10'b0000000001, locator0, alpha284_0_x_locator0);
  gfmult gfm_alpha284_1_x_locator1(10'b1011101010, locator1, alpha284_1_x_locator1);
  gfmult gfm_alpha284_2_x_locator2(10'b0111101011, locator2, alpha284_2_x_locator2);
  gfmult gfm_alpha284_3_x_locator3(10'b1010101101, locator3, alpha284_3_x_locator3);
  gfmult gfm_alpha285_0_x_locator0(10'b0000000001, locator0, alpha285_0_x_locator0);
  gfmult gfm_alpha285_1_x_locator1(10'b0101110101, locator1, alpha285_1_x_locator1);
  gfmult gfm_alpha285_2_x_locator2(10'b1101111100, locator2, alpha285_2_x_locator2);
  gfmult gfm_alpha285_3_x_locator3(10'b1011010000, locator3, alpha285_3_x_locator3);
  gfmult gfm_alpha286_0_x_locator0(10'b0000000001, locator0, alpha286_0_x_locator0);
  gfmult gfm_alpha286_1_x_locator1(10'b1010111110, locator1, alpha286_1_x_locator1);
  gfmult gfm_alpha286_2_x_locator2(10'b0011011111, locator2, alpha286_2_x_locator2);
  gfmult gfm_alpha286_3_x_locator3(10'b0001011010, locator3, alpha286_3_x_locator3);
  gfmult gfm_alpha287_0_x_locator0(10'b0000000001, locator0, alpha287_0_x_locator0);
  gfmult gfm_alpha287_1_x_locator1(10'b0101011111, locator1, alpha287_1_x_locator1);
  gfmult gfm_alpha287_2_x_locator2(10'b1100110001, locator2, alpha287_2_x_locator2);
  gfmult gfm_alpha287_3_x_locator3(10'b0100001001, locator3, alpha287_3_x_locator3);
  gfmult gfm_alpha288_0_x_locator0(10'b0000000001, locator0, alpha288_0_x_locator0);
  gfmult gfm_alpha288_1_x_locator1(10'b1010101011, locator1, alpha288_1_x_locator1);
  gfmult gfm_alpha288_2_x_locator2(10'b0111001110, locator2, alpha288_2_x_locator2);
  gfmult gfm_alpha288_3_x_locator3(10'b0010100000, locator3, alpha288_3_x_locator3);
  gfmult gfm_alpha289_0_x_locator0(10'b0000000001, locator0, alpha289_0_x_locator0);
  gfmult gfm_alpha289_1_x_locator1(10'b1101010001, locator1, alpha289_1_x_locator1);
  gfmult gfm_alpha289_2_x_locator2(10'b1001110111, locator2, alpha289_2_x_locator2);
  gfmult gfm_alpha289_3_x_locator3(10'b0000010100, locator3, alpha289_3_x_locator3);
  gfmult gfm_alpha290_0_x_locator0(10'b0000000001, locator0, alpha290_0_x_locator0);
  gfmult gfm_alpha290_1_x_locator1(10'b1110101100, locator1, alpha290_1_x_locator1);
  gfmult gfm_alpha290_2_x_locator2(10'b1110011011, locator2, alpha290_2_x_locator2);
  gfmult gfm_alpha290_3_x_locator3(10'b1000000110, locator3, alpha290_3_x_locator3);
  gfmult gfm_alpha291_0_x_locator0(10'b0000000001, locator0, alpha291_0_x_locator0);
  gfmult gfm_alpha291_1_x_locator1(10'b0111010110, locator1, alpha291_1_x_locator1);
  gfmult gfm_alpha291_2_x_locator2(10'b1111100000, locator2, alpha291_2_x_locator2);
  gfmult gfm_alpha291_3_x_locator3(10'b1101000110, locator3, alpha291_3_x_locator3);
  gfmult gfm_alpha292_0_x_locator0(10'b0000000001, locator0, alpha292_0_x_locator0);
  gfmult gfm_alpha292_1_x_locator1(10'b0011101011, locator1, alpha292_1_x_locator1);
  gfmult gfm_alpha292_2_x_locator2(10'b0011111000, locator2, alpha292_2_x_locator2);
  gfmult gfm_alpha292_3_x_locator3(10'b1101101110, locator3, alpha292_3_x_locator3);
  gfmult gfm_alpha293_0_x_locator0(10'b0000000001, locator0, alpha293_0_x_locator0);
  gfmult gfm_alpha293_1_x_locator1(10'b1001110001, locator1, alpha293_1_x_locator1);
  gfmult gfm_alpha293_2_x_locator2(10'b0000111110, locator2, alpha293_2_x_locator2);
  gfmult gfm_alpha293_3_x_locator3(10'b1101101011, locator3, alpha293_3_x_locator3);
  gfmult gfm_alpha294_0_x_locator0(10'b0000000001, locator0, alpha294_0_x_locator0);
  gfmult gfm_alpha294_1_x_locator1(10'b1100111100, locator1, alpha294_1_x_locator1);
  gfmult gfm_alpha294_2_x_locator2(10'b1000001011, locator2, alpha294_2_x_locator2);
  gfmult gfm_alpha294_3_x_locator3(10'b0111101110, locator3, alpha294_3_x_locator3);
  gfmult gfm_alpha295_0_x_locator0(10'b0000000001, locator0, alpha295_0_x_locator0);
  gfmult gfm_alpha295_1_x_locator1(10'b0110011110, locator1, alpha295_1_x_locator1);
  gfmult gfm_alpha295_2_x_locator2(10'b1110000100, locator2, alpha295_2_x_locator2);
  gfmult gfm_alpha295_3_x_locator3(10'b1100111011, locator3, alpha295_3_x_locator3);
  gfmult gfm_alpha296_0_x_locator0(10'b0000000001, locator0, alpha296_0_x_locator0);
  gfmult gfm_alpha296_1_x_locator1(10'b0011001111, locator1, alpha296_1_x_locator1);
  gfmult gfm_alpha296_2_x_locator2(10'b0011100001, locator2, alpha296_2_x_locator2);
  gfmult gfm_alpha296_3_x_locator3(10'b0111100100, locator3, alpha296_3_x_locator3);
  gfmult gfm_alpha297_0_x_locator0(10'b0000000001, locator0, alpha297_0_x_locator0);
  gfmult gfm_alpha297_1_x_locator1(10'b1001100011, locator1, alpha297_1_x_locator1);
  gfmult gfm_alpha297_2_x_locator2(10'b0100111010, locator2, alpha297_2_x_locator2);
  gfmult gfm_alpha297_3_x_locator3(10'b1000111000, locator3, alpha297_3_x_locator3);
  gfmult gfm_alpha298_0_x_locator0(10'b0000000001, locator0, alpha298_0_x_locator0);
  gfmult gfm_alpha298_1_x_locator1(10'b1100110101, locator1, alpha298_1_x_locator1);
  gfmult gfm_alpha298_2_x_locator2(10'b1001001010, locator2, alpha298_2_x_locator2);
  gfmult gfm_alpha298_3_x_locator3(10'b0001000111, locator3, alpha298_3_x_locator3);
  gfmult gfm_alpha299_0_x_locator0(10'b0000000001, locator0, alpha299_0_x_locator0);
  gfmult gfm_alpha299_1_x_locator1(10'b1110011110, locator1, alpha299_1_x_locator1);
  gfmult gfm_alpha299_2_x_locator2(10'b1010010110, locator2, alpha299_2_x_locator2);
  gfmult gfm_alpha299_3_x_locator3(10'b1110001111, locator3, alpha299_3_x_locator3);
  gfmult gfm_alpha300_0_x_locator0(10'b0000000001, locator0, alpha300_0_x_locator0);
  gfmult gfm_alpha300_1_x_locator1(10'b0111001111, locator1, alpha300_1_x_locator1);
  gfmult gfm_alpha300_2_x_locator2(10'b1010100001, locator2, alpha300_2_x_locator2);
  gfmult gfm_alpha300_3_x_locator3(10'b1111110110, locator3, alpha300_3_x_locator3);
  gfmult gfm_alpha301_0_x_locator0(10'b0000000001, locator0, alpha301_0_x_locator0);
  gfmult gfm_alpha301_1_x_locator1(10'b1011100011, locator1, alpha301_1_x_locator1);
  gfmult gfm_alpha301_2_x_locator2(10'b0110101010, locator2, alpha301_2_x_locator2);
  gfmult gfm_alpha301_3_x_locator3(10'b1101111000, locator3, alpha301_3_x_locator3);
  gfmult gfm_alpha302_0_x_locator0(10'b0000000001, locator0, alpha302_0_x_locator0);
  gfmult gfm_alpha302_1_x_locator1(10'b1101110101, locator1, alpha302_1_x_locator1);
  gfmult gfm_alpha302_2_x_locator2(10'b1001101110, locator2, alpha302_2_x_locator2);
  gfmult gfm_alpha302_3_x_locator3(10'b0001101111, locator3, alpha302_3_x_locator3);
  gfmult gfm_alpha303_0_x_locator0(10'b0000000001, locator0, alpha303_0_x_locator0);
  gfmult gfm_alpha303_1_x_locator1(10'b1110111110, locator1, alpha303_1_x_locator1);
  gfmult gfm_alpha303_2_x_locator2(10'b1010011111, locator2, alpha303_2_x_locator2);
  gfmult gfm_alpha303_3_x_locator3(10'b1110001010, locator3, alpha303_3_x_locator3);
  gfmult gfm_alpha304_0_x_locator0(10'b0000000001, locator0, alpha304_0_x_locator0);
  gfmult gfm_alpha304_1_x_locator1(10'b0111011111, locator1, alpha304_1_x_locator1);
  gfmult gfm_alpha304_2_x_locator2(10'b1110100001, locator2, alpha304_2_x_locator2);
  gfmult gfm_alpha304_3_x_locator3(10'b0101110011, locator3, alpha304_3_x_locator3);
  gfmult gfm_alpha305_0_x_locator0(10'b0000000001, locator0, alpha305_0_x_locator0);
  gfmult gfm_alpha305_1_x_locator1(10'b1011101011, locator1, alpha305_1_x_locator1);
  gfmult gfm_alpha305_2_x_locator2(10'b0111101010, locator2, alpha305_2_x_locator2);
  gfmult gfm_alpha305_3_x_locator3(10'b0110101101, locator3, alpha305_3_x_locator3);
  gfmult gfm_alpha306_0_x_locator0(10'b0000000001, locator0, alpha306_0_x_locator0);
  gfmult gfm_alpha306_1_x_locator1(10'b1101110001, locator1, alpha306_1_x_locator1);
  gfmult gfm_alpha306_2_x_locator2(10'b1001111110, locator2, alpha306_2_x_locator2);
  gfmult gfm_alpha306_3_x_locator3(10'b1010110000, locator3, alpha306_3_x_locator3);
  gfmult gfm_alpha307_0_x_locator0(10'b0000000001, locator0, alpha307_0_x_locator0);
  gfmult gfm_alpha307_1_x_locator1(10'b1110111100, locator1, alpha307_1_x_locator1);
  gfmult gfm_alpha307_2_x_locator2(10'b1010011011, locator2, alpha307_2_x_locator2);
  gfmult gfm_alpha307_3_x_locator3(10'b0001010110, locator3, alpha307_3_x_locator3);
  gfmult gfm_alpha308_0_x_locator0(10'b0000000001, locator0, alpha308_0_x_locator0);
  gfmult gfm_alpha308_1_x_locator1(10'b0111011110, locator1, alpha308_1_x_locator1);
  gfmult gfm_alpha308_2_x_locator2(10'b1110100000, locator2, alpha308_2_x_locator2);
  gfmult gfm_alpha308_3_x_locator3(10'b1100001100, locator3, alpha308_3_x_locator3);
  gfmult gfm_alpha309_0_x_locator0(10'b0000000001, locator0, alpha309_0_x_locator0);
  gfmult gfm_alpha309_1_x_locator1(10'b0011101111, locator1, alpha309_1_x_locator1);
  gfmult gfm_alpha309_2_x_locator2(10'b0011101000, locator2, alpha309_2_x_locator2);
  gfmult gfm_alpha309_3_x_locator3(10'b1001100101, locator3, alpha309_3_x_locator3);
  gfmult gfm_alpha310_0_x_locator0(10'b0000000001, locator0, alpha310_0_x_locator0);
  gfmult gfm_alpha310_1_x_locator1(10'b1001110011, locator1, alpha310_1_x_locator1);
  gfmult gfm_alpha310_2_x_locator2(10'b0000111010, locator2, alpha310_2_x_locator2);
  gfmult gfm_alpha310_3_x_locator3(10'b1011001001, locator3, alpha310_3_x_locator3);
  gfmult gfm_alpha311_0_x_locator0(10'b0000000001, locator0, alpha311_0_x_locator0);
  gfmult gfm_alpha311_1_x_locator1(10'b1100111101, locator1, alpha311_1_x_locator1);
  gfmult gfm_alpha311_2_x_locator2(10'b1000001010, locator2, alpha311_2_x_locator2);
  gfmult gfm_alpha311_3_x_locator3(10'b0011011000, locator3, alpha311_3_x_locator3);
  gfmult gfm_alpha312_0_x_locator0(10'b0000000001, locator0, alpha312_0_x_locator0);
  gfmult gfm_alpha312_1_x_locator1(10'b1110011010, locator1, alpha312_1_x_locator1);
  gfmult gfm_alpha312_2_x_locator2(10'b1010000110, locator2, alpha312_2_x_locator2);
  gfmult gfm_alpha312_3_x_locator3(10'b0000011011, locator3, alpha312_3_x_locator3);
  gfmult gfm_alpha313_0_x_locator0(10'b0000000001, locator0, alpha313_0_x_locator0);
  gfmult gfm_alpha313_1_x_locator1(10'b0111001101, locator1, alpha313_1_x_locator1);
  gfmult gfm_alpha313_2_x_locator2(10'b1010100101, locator2, alpha313_2_x_locator2);
  gfmult gfm_alpha313_3_x_locator3(10'b0110000000, locator3, alpha313_3_x_locator3);
  gfmult gfm_alpha314_0_x_locator0(10'b0000000001, locator0, alpha314_0_x_locator0);
  gfmult gfm_alpha314_1_x_locator1(10'b1011100010, locator1, alpha314_1_x_locator1);
  gfmult gfm_alpha314_2_x_locator2(10'b0110101011, locator2, alpha314_2_x_locator2);
  gfmult gfm_alpha314_3_x_locator3(10'b0000110000, locator3, alpha314_3_x_locator3);
  gfmult gfm_alpha315_0_x_locator0(10'b0000000001, locator0, alpha315_0_x_locator0);
  gfmult gfm_alpha315_1_x_locator1(10'b0101110001, locator1, alpha315_1_x_locator1);
  gfmult gfm_alpha315_2_x_locator2(10'b1101101100, locator2, alpha315_2_x_locator2);
  gfmult gfm_alpha315_3_x_locator3(10'b0000000110, locator3, alpha315_3_x_locator3);
  gfmult gfm_alpha316_0_x_locator0(10'b0000000001, locator0, alpha316_0_x_locator0);
  gfmult gfm_alpha316_1_x_locator1(10'b1010111100, locator1, alpha316_1_x_locator1);
  gfmult gfm_alpha316_2_x_locator2(10'b0011011011, locator2, alpha316_2_x_locator2);
  gfmult gfm_alpha316_3_x_locator3(10'b1100000110, locator3, alpha316_3_x_locator3);
  gfmult gfm_alpha317_0_x_locator0(10'b0000000001, locator0, alpha317_0_x_locator0);
  gfmult gfm_alpha317_1_x_locator1(10'b0101011110, locator1, alpha317_1_x_locator1);
  gfmult gfm_alpha317_2_x_locator2(10'b1100110000, locator2, alpha317_2_x_locator2);
  gfmult gfm_alpha317_3_x_locator3(10'b1101100110, locator3, alpha317_3_x_locator3);
  gfmult gfm_alpha318_0_x_locator0(10'b0000000001, locator0, alpha318_0_x_locator0);
  gfmult gfm_alpha318_1_x_locator1(10'b0010101111, locator1, alpha318_1_x_locator1);
  gfmult gfm_alpha318_2_x_locator2(10'b0011001100, locator2, alpha318_2_x_locator2);
  gfmult gfm_alpha318_3_x_locator3(10'b1101101010, locator3, alpha318_3_x_locator3);
  gfmult gfm_alpha319_0_x_locator0(10'b0000000001, locator0, alpha319_0_x_locator0);
  gfmult gfm_alpha319_1_x_locator1(10'b1001010011, locator1, alpha319_1_x_locator1);
  gfmult gfm_alpha319_2_x_locator2(10'b0000110011, locator2, alpha319_2_x_locator2);
  gfmult gfm_alpha319_3_x_locator3(10'b0101101111, locator3, alpha319_3_x_locator3);
  gfmult gfm_alpha320_0_x_locator0(10'b0000000001, locator0, alpha320_0_x_locator0);
  gfmult gfm_alpha320_1_x_locator1(10'b1100101101, locator1, alpha320_1_x_locator1);
  gfmult gfm_alpha320_2_x_locator2(10'b1100001010, locator2, alpha320_2_x_locator2);
  gfmult gfm_alpha320_3_x_locator3(10'b1110101010, locator3, alpha320_3_x_locator3);
  gfmult gfm_alpha321_0_x_locator0(10'b0000000001, locator0, alpha321_0_x_locator0);
  gfmult gfm_alpha321_1_x_locator1(10'b1110010010, locator1, alpha321_1_x_locator1);
  gfmult gfm_alpha321_2_x_locator2(10'b1011000110, locator2, alpha321_2_x_locator2);
  gfmult gfm_alpha321_3_x_locator3(10'b0101110111, locator3, alpha321_3_x_locator3);
  gfmult gfm_alpha322_0_x_locator0(10'b0000000001, locator0, alpha322_0_x_locator0);
  gfmult gfm_alpha322_1_x_locator1(10'b0111001001, locator1, alpha322_1_x_locator1);
  gfmult gfm_alpha322_2_x_locator2(10'b1010110101, locator2, alpha322_2_x_locator2);
  gfmult gfm_alpha322_3_x_locator3(10'b1110101001, locator3, alpha322_3_x_locator3);
  gfmult gfm_alpha323_0_x_locator0(10'b0000000001, locator0, alpha323_0_x_locator0);
  gfmult gfm_alpha323_1_x_locator1(10'b1011100000, locator1, alpha323_1_x_locator1);
  gfmult gfm_alpha323_2_x_locator2(10'b0110101111, locator2, alpha323_2_x_locator2);
  gfmult gfm_alpha323_3_x_locator3(10'b0011110100, locator3, alpha323_3_x_locator3);
  gfmult gfm_alpha324_0_x_locator0(10'b0000000001, locator0, alpha324_0_x_locator0);
  gfmult gfm_alpha324_1_x_locator1(10'b0101110000, locator1, alpha324_1_x_locator1);
  gfmult gfm_alpha324_2_x_locator2(10'b1101101101, locator2, alpha324_2_x_locator2);
  gfmult gfm_alpha324_3_x_locator3(10'b1000011010, locator3, alpha324_3_x_locator3);
  gfmult gfm_alpha325_0_x_locator0(10'b0000000001, locator0, alpha325_0_x_locator0);
  gfmult gfm_alpha325_1_x_locator1(10'b0010111000, locator1, alpha325_1_x_locator1);
  gfmult gfm_alpha325_2_x_locator2(10'b0111011001, locator2, alpha325_2_x_locator2);
  gfmult gfm_alpha325_3_x_locator3(10'b0101000001, locator3, alpha325_3_x_locator3);
  gfmult gfm_alpha326_0_x_locator0(10'b0000000001, locator0, alpha326_0_x_locator0);
  gfmult gfm_alpha326_1_x_locator1(10'b0001011100, locator1, alpha326_1_x_locator1);
  gfmult gfm_alpha326_2_x_locator2(10'b0101110100, locator2, alpha326_2_x_locator2);
  gfmult gfm_alpha326_3_x_locator3(10'b0010101001, locator3, alpha326_3_x_locator3);
  gfmult gfm_alpha327_0_x_locator0(10'b0000000001, locator0, alpha327_0_x_locator0);
  gfmult gfm_alpha327_1_x_locator1(10'b0000101110, locator1, alpha327_1_x_locator1);
  gfmult gfm_alpha327_2_x_locator2(10'b0001011101, locator2, alpha327_2_x_locator2);
  gfmult gfm_alpha327_3_x_locator3(10'b0010010100, locator3, alpha327_3_x_locator3);
  gfmult gfm_alpha328_0_x_locator0(10'b0000000001, locator0, alpha328_0_x_locator0);
  gfmult gfm_alpha328_1_x_locator1(10'b0000010111, locator1, alpha328_1_x_locator1);
  gfmult gfm_alpha328_2_x_locator2(10'b0100010101, locator2, alpha328_2_x_locator2);
  gfmult gfm_alpha328_3_x_locator3(10'b1000010110, locator3, alpha328_3_x_locator3);
  gfmult gfm_alpha329_0_x_locator0(10'b0000000001, locator0, alpha329_0_x_locator0);
  gfmult gfm_alpha329_1_x_locator1(10'b1000001111, locator1, alpha329_1_x_locator1);
  gfmult gfm_alpha329_2_x_locator2(10'b0101000111, locator2, alpha329_2_x_locator2);
  gfmult gfm_alpha329_3_x_locator3(10'b1101000100, locator3, alpha329_3_x_locator3);
  gfmult gfm_alpha330_0_x_locator0(10'b0000000001, locator0, alpha330_0_x_locator0);
  gfmult gfm_alpha330_1_x_locator1(10'b1100000011, locator1, alpha330_1_x_locator1);
  gfmult gfm_alpha330_2_x_locator2(10'b1101010111, locator2, alpha330_2_x_locator2);
  gfmult gfm_alpha330_3_x_locator3(10'b1001101100, locator3, alpha330_3_x_locator3);
  gfmult gfm_alpha331_0_x_locator0(10'b0000000001, locator0, alpha331_0_x_locator0);
  gfmult gfm_alpha331_1_x_locator1(10'b1110000101, locator1, alpha331_1_x_locator1);
  gfmult gfm_alpha331_2_x_locator2(10'b1111010011, locator2, alpha331_2_x_locator2);
  gfmult gfm_alpha331_3_x_locator3(10'b1001001001, locator3, alpha331_3_x_locator3);
  gfmult gfm_alpha332_0_x_locator0(10'b0000000001, locator0, alpha332_0_x_locator0);
  gfmult gfm_alpha332_1_x_locator1(10'b1111000110, locator1, alpha332_1_x_locator1);
  gfmult gfm_alpha332_2_x_locator2(10'b1111110010, locator2, alpha332_2_x_locator2);
  gfmult gfm_alpha332_3_x_locator3(10'b0011001000, locator3, alpha332_3_x_locator3);
  gfmult gfm_alpha333_0_x_locator0(10'b0000000001, locator0, alpha333_0_x_locator0);
  gfmult gfm_alpha333_1_x_locator1(10'b0111100011, locator1, alpha333_1_x_locator1);
  gfmult gfm_alpha333_2_x_locator2(10'b1011111000, locator2, alpha333_2_x_locator2);
  gfmult gfm_alpha333_3_x_locator3(10'b0000011001, locator3, alpha333_3_x_locator3);
  gfmult gfm_alpha334_0_x_locator0(10'b0000000001, locator0, alpha334_0_x_locator0);
  gfmult gfm_alpha334_1_x_locator1(10'b1011110101, locator1, alpha334_1_x_locator1);
  gfmult gfm_alpha334_2_x_locator2(10'b0010111110, locator2, alpha334_2_x_locator2);
  gfmult gfm_alpha334_3_x_locator3(10'b0010000010, locator3, alpha334_3_x_locator3);
  gfmult gfm_alpha335_0_x_locator0(10'b0000000001, locator0, alpha335_0_x_locator0);
  gfmult gfm_alpha335_1_x_locator1(10'b1101111110, locator1, alpha335_1_x_locator1);
  gfmult gfm_alpha335_2_x_locator2(10'b1000101011, locator2, alpha335_2_x_locator2);
  gfmult gfm_alpha335_3_x_locator3(10'b0100010010, locator3, alpha335_3_x_locator3);
  gfmult gfm_alpha336_0_x_locator0(10'b0000000001, locator0, alpha336_0_x_locator0);
  gfmult gfm_alpha336_1_x_locator1(10'b0110111111, locator1, alpha336_1_x_locator1);
  gfmult gfm_alpha336_2_x_locator2(10'b1110001100, locator2, alpha336_2_x_locator2);
  gfmult gfm_alpha336_3_x_locator3(10'b0100100000, locator3, alpha336_3_x_locator3);
  gfmult gfm_alpha337_0_x_locator0(10'b0000000001, locator0, alpha337_0_x_locator0);
  gfmult gfm_alpha337_1_x_locator1(10'b1011011011, locator1, alpha337_1_x_locator1);
  gfmult gfm_alpha337_2_x_locator2(10'b0011100011, locator2, alpha337_2_x_locator2);
  gfmult gfm_alpha337_3_x_locator3(10'b0000100100, locator3, alpha337_3_x_locator3);
  gfmult gfm_alpha338_0_x_locator0(10'b0000000001, locator0, alpha338_0_x_locator0);
  gfmult gfm_alpha338_1_x_locator1(10'b1101101001, locator1, alpha338_1_x_locator1);
  gfmult gfm_alpha338_2_x_locator2(10'b1100111110, locator2, alpha338_2_x_locator2);
  gfmult gfm_alpha338_3_x_locator3(10'b1000000000, locator3, alpha338_3_x_locator3);
  gfmult gfm_alpha339_0_x_locator0(10'b0000000001, locator0, alpha339_0_x_locator0);
  gfmult gfm_alpha339_1_x_locator1(10'b1110110000, locator1, alpha339_1_x_locator1);
  gfmult gfm_alpha339_2_x_locator2(10'b1011001011, locator2, alpha339_2_x_locator2);
  gfmult gfm_alpha339_3_x_locator3(10'b0001000000, locator3, alpha339_3_x_locator3);
  gfmult gfm_alpha340_0_x_locator0(10'b0000000001, locator0, alpha340_0_x_locator0);
  gfmult gfm_alpha340_1_x_locator1(10'b0111011000, locator1, alpha340_1_x_locator1);
  gfmult gfm_alpha340_2_x_locator2(10'b1110110100, locator2, alpha340_2_x_locator2);
  gfmult gfm_alpha340_3_x_locator3(10'b0000001000, locator3, alpha340_3_x_locator3);
  gfmult gfm_alpha341_0_x_locator0(10'b0000000001, locator0, alpha341_0_x_locator0);
  gfmult gfm_alpha341_1_x_locator1(10'b0011101100, locator1, alpha341_1_x_locator1);
  gfmult gfm_alpha341_2_x_locator2(10'b0011101101, locator2, alpha341_2_x_locator2);
  gfmult gfm_alpha341_3_x_locator3(10'b0000000001, locator3, alpha341_3_x_locator3);
  gfmult gfm_alpha342_0_x_locator0(10'b0000000001, locator0, alpha342_0_x_locator0);
  gfmult gfm_alpha342_1_x_locator1(10'b0001110110, locator1, alpha342_1_x_locator1);
  gfmult gfm_alpha342_2_x_locator2(10'b0100111001, locator2, alpha342_2_x_locator2);
  gfmult gfm_alpha342_3_x_locator3(10'b0010000001, locator3, alpha342_3_x_locator3);
  gfmult gfm_alpha343_0_x_locator0(10'b0000000001, locator0, alpha343_0_x_locator0);
  gfmult gfm_alpha343_1_x_locator1(10'b0000111011, locator1, alpha343_1_x_locator1);
  gfmult gfm_alpha343_2_x_locator2(10'b0101001100, locator2, alpha343_2_x_locator2);
  gfmult gfm_alpha343_3_x_locator3(10'b0010010001, locator3, alpha343_3_x_locator3);
  gfmult gfm_alpha344_0_x_locator0(10'b0000000001, locator0, alpha344_0_x_locator0);
  gfmult gfm_alpha344_1_x_locator1(10'b1000011001, locator1, alpha344_1_x_locator1);
  gfmult gfm_alpha344_2_x_locator2(10'b0001010011, locator2, alpha344_2_x_locator2);
  gfmult gfm_alpha344_3_x_locator3(10'b0010010011, locator3, alpha344_3_x_locator3);
  gfmult gfm_alpha345_0_x_locator0(10'b0000000001, locator0, alpha345_0_x_locator0);
  gfmult gfm_alpha345_1_x_locator1(10'b1100001000, locator1, alpha345_1_x_locator1);
  gfmult gfm_alpha345_2_x_locator2(10'b1100010010, locator2, alpha345_2_x_locator2);
  gfmult gfm_alpha345_3_x_locator3(10'b0110010001, locator3, alpha345_3_x_locator3);
  gfmult gfm_alpha346_0_x_locator0(10'b0000000001, locator0, alpha346_0_x_locator0);
  gfmult gfm_alpha346_1_x_locator1(10'b0110000100, locator1, alpha346_1_x_locator1);
  gfmult gfm_alpha346_2_x_locator2(10'b1011000000, locator2, alpha346_2_x_locator2);
  gfmult gfm_alpha346_3_x_locator3(10'b0010110011, locator3, alpha346_3_x_locator3);
  gfmult gfm_alpha347_0_x_locator0(10'b0000000001, locator0, alpha347_0_x_locator0);
  gfmult gfm_alpha347_1_x_locator1(10'b0011000010, locator1, alpha347_1_x_locator1);
  gfmult gfm_alpha347_2_x_locator2(10'b0010110000, locator2, alpha347_2_x_locator2);
  gfmult gfm_alpha347_3_x_locator3(10'b0110010101, locator3, alpha347_3_x_locator3);
  gfmult gfm_alpha348_0_x_locator0(10'b0000000001, locator0, alpha348_0_x_locator0);
  gfmult gfm_alpha348_1_x_locator1(10'b0001100001, locator1, alpha348_1_x_locator1);
  gfmult gfm_alpha348_2_x_locator2(10'b0000101100, locator2, alpha348_2_x_locator2);
  gfmult gfm_alpha348_3_x_locator3(10'b1010110111, locator3, alpha348_3_x_locator3);
  gfmult gfm_alpha349_0_x_locator0(10'b0000000001, locator0, alpha349_0_x_locator0);
  gfmult gfm_alpha349_1_x_locator1(10'b1000110100, locator1, alpha349_1_x_locator1);
  gfmult gfm_alpha349_2_x_locator2(10'b0000001011, locator2, alpha349_2_x_locator2);
  gfmult gfm_alpha349_3_x_locator3(10'b1111010001, locator3, alpha349_3_x_locator3);
  gfmult gfm_alpha350_0_x_locator0(10'b0000000001, locator0, alpha350_0_x_locator0);
  gfmult gfm_alpha350_1_x_locator1(10'b0100011010, locator1, alpha350_1_x_locator1);
  gfmult gfm_alpha350_2_x_locator2(10'b1100000100, locator2, alpha350_2_x_locator2);
  gfmult gfm_alpha350_3_x_locator3(10'b0011111011, locator3, alpha350_3_x_locator3);
  gfmult gfm_alpha351_0_x_locator0(10'b0000000001, locator0, alpha351_0_x_locator0);
  gfmult gfm_alpha351_1_x_locator1(10'b0010001101, locator1, alpha351_1_x_locator1);
  gfmult gfm_alpha351_2_x_locator2(10'b0011000001, locator2, alpha351_2_x_locator2);
  gfmult gfm_alpha351_3_x_locator3(10'b0110011100, locator3, alpha351_3_x_locator3);
  gfmult gfm_alpha352_0_x_locator0(10'b0000000001, locator0, alpha352_0_x_locator0);
  gfmult gfm_alpha352_1_x_locator1(10'b1001000010, locator1, alpha352_1_x_locator1);
  gfmult gfm_alpha352_2_x_locator2(10'b0100110010, locator2, alpha352_2_x_locator2);
  gfmult gfm_alpha352_3_x_locator3(10'b1000110111, locator3, alpha352_3_x_locator3);
  gfmult gfm_alpha353_0_x_locator0(10'b0000000001, locator0, alpha353_0_x_locator0);
  gfmult gfm_alpha353_1_x_locator1(10'b0100100001, locator1, alpha353_1_x_locator1);
  gfmult gfm_alpha353_2_x_locator2(10'b1001001000, locator2, alpha353_2_x_locator2);
  gfmult gfm_alpha353_3_x_locator3(10'b1111000001, locator3, alpha353_3_x_locator3);
  gfmult gfm_alpha354_0_x_locator0(10'b0000000001, locator0, alpha354_0_x_locator0);
  gfmult gfm_alpha354_1_x_locator1(10'b1010010100, locator1, alpha354_1_x_locator1);
  gfmult gfm_alpha354_2_x_locator2(10'b0010010010, locator2, alpha354_2_x_locator2);
  gfmult gfm_alpha354_3_x_locator3(10'b0011111001, locator3, alpha354_3_x_locator3);
  gfmult gfm_alpha355_0_x_locator0(10'b0000000001, locator0, alpha355_0_x_locator0);
  gfmult gfm_alpha355_1_x_locator1(10'b0101001010, locator1, alpha355_1_x_locator1);
  gfmult gfm_alpha355_2_x_locator2(10'b1000100000, locator2, alpha355_2_x_locator2);
  gfmult gfm_alpha355_3_x_locator3(10'b0010011110, locator3, alpha355_3_x_locator3);
  gfmult gfm_alpha356_0_x_locator0(10'b0000000001, locator0, alpha356_0_x_locator0);
  gfmult gfm_alpha356_1_x_locator1(10'b0010100101, locator1, alpha356_1_x_locator1);
  gfmult gfm_alpha356_2_x_locator2(10'b0010001000, locator2, alpha356_2_x_locator2);
  gfmult gfm_alpha356_3_x_locator3(10'b1100010101, locator3, alpha356_3_x_locator3);
  gfmult gfm_alpha357_0_x_locator0(10'b0000000001, locator0, alpha357_0_x_locator0);
  gfmult gfm_alpha357_1_x_locator1(10'b1001010110, locator1, alpha357_1_x_locator1);
  gfmult gfm_alpha357_2_x_locator2(10'b0000100010, locator2, alpha357_2_x_locator2);
  gfmult gfm_alpha357_3_x_locator3(10'b1011100111, locator3, alpha357_3_x_locator3);
  gfmult gfm_alpha358_0_x_locator0(10'b0000000001, locator0, alpha358_0_x_locator0);
  gfmult gfm_alpha358_1_x_locator1(10'b0100101011, locator1, alpha358_1_x_locator1);
  gfmult gfm_alpha358_2_x_locator2(10'b1000001100, locator2, alpha358_2_x_locator2);
  gfmult gfm_alpha358_3_x_locator3(10'b1111011011, locator3, alpha358_3_x_locator3);
  gfmult gfm_alpha359_0_x_locator0(10'b0000000001, locator0, alpha359_0_x_locator0);
  gfmult gfm_alpha359_1_x_locator1(10'b1010010001, locator1, alpha359_1_x_locator1);
  gfmult gfm_alpha359_2_x_locator2(10'b0010000011, locator2, alpha359_2_x_locator2);
  gfmult gfm_alpha359_3_x_locator3(10'b0111111000, locator3, alpha359_3_x_locator3);
  gfmult gfm_alpha360_0_x_locator0(10'b0000000001, locator0, alpha360_0_x_locator0);
  gfmult gfm_alpha360_1_x_locator1(10'b1101001100, locator1, alpha360_1_x_locator1);
  gfmult gfm_alpha360_2_x_locator2(10'b1100100110, locator2, alpha360_2_x_locator2);
  gfmult gfm_alpha360_3_x_locator3(10'b0000111111, locator3, alpha360_3_x_locator3);
  gfmult gfm_alpha361_0_x_locator0(10'b0000000001, locator0, alpha361_0_x_locator0);
  gfmult gfm_alpha361_1_x_locator1(10'b0110100110, locator1, alpha361_1_x_locator1);
  gfmult gfm_alpha361_2_x_locator2(10'b1011001101, locator2, alpha361_2_x_locator2);
  gfmult gfm_alpha361_3_x_locator3(10'b1110000000, locator3, alpha361_3_x_locator3);
  gfmult gfm_alpha362_0_x_locator0(10'b0000000001, locator0, alpha362_0_x_locator0);
  gfmult gfm_alpha362_1_x_locator1(10'b0011010011, locator1, alpha362_1_x_locator1);
  gfmult gfm_alpha362_2_x_locator2(10'b0110110001, locator2, alpha362_2_x_locator2);
  gfmult gfm_alpha362_3_x_locator3(10'b0001110000, locator3, alpha362_3_x_locator3);
  gfmult gfm_alpha363_0_x_locator0(10'b0000000001, locator0, alpha363_0_x_locator0);
  gfmult gfm_alpha363_1_x_locator1(10'b1001101101, locator1, alpha363_1_x_locator1);
  gfmult gfm_alpha363_2_x_locator2(10'b0101101110, locator2, alpha363_2_x_locator2);
  gfmult gfm_alpha363_3_x_locator3(10'b0000001110, locator3, alpha363_3_x_locator3);
  gfmult gfm_alpha364_0_x_locator0(10'b0000000001, locator0, alpha364_0_x_locator0);
  gfmult gfm_alpha364_1_x_locator1(10'b1100110010, locator1, alpha364_1_x_locator1);
  gfmult gfm_alpha364_2_x_locator2(10'b1001011111, locator2, alpha364_2_x_locator2);
  gfmult gfm_alpha364_3_x_locator3(10'b1100000111, locator3, alpha364_3_x_locator3);
  gfmult gfm_alpha365_0_x_locator0(10'b0000000001, locator0, alpha365_0_x_locator0);
  gfmult gfm_alpha365_1_x_locator1(10'b0110011001, locator1, alpha365_1_x_locator1);
  gfmult gfm_alpha365_2_x_locator2(10'b1110010001, locator2, alpha365_2_x_locator2);
  gfmult gfm_alpha365_3_x_locator3(10'b1111100111, locator3, alpha365_3_x_locator3);
  gfmult gfm_alpha366_0_x_locator0(10'b0000000001, locator0, alpha366_0_x_locator0);
  gfmult gfm_alpha366_1_x_locator1(10'b1011001000, locator1, alpha366_1_x_locator1);
  gfmult gfm_alpha366_2_x_locator2(10'b0111100110, locator2, alpha366_2_x_locator2);
  gfmult gfm_alpha366_3_x_locator3(10'b1111111011, locator3, alpha366_3_x_locator3);
  gfmult gfm_alpha367_0_x_locator0(10'b0000000001, locator0, alpha367_0_x_locator0);
  gfmult gfm_alpha367_1_x_locator1(10'b0101100100, locator1, alpha367_1_x_locator1);
  gfmult gfm_alpha367_2_x_locator2(10'b1001111101, locator2, alpha367_2_x_locator2);
  gfmult gfm_alpha367_3_x_locator3(10'b0111111100, locator3, alpha367_3_x_locator3);
  gfmult gfm_alpha368_0_x_locator0(10'b0000000001, locator0, alpha368_0_x_locator0);
  gfmult gfm_alpha368_1_x_locator1(10'b0010110010, locator1, alpha368_1_x_locator1);
  gfmult gfm_alpha368_2_x_locator2(10'b0110011101, locator2, alpha368_2_x_locator2);
  gfmult gfm_alpha368_3_x_locator3(10'b1000111011, locator3, alpha368_3_x_locator3);
  gfmult gfm_alpha369_0_x_locator0(10'b0000000001, locator0, alpha369_0_x_locator0);
  gfmult gfm_alpha369_1_x_locator1(10'b0001011001, locator1, alpha369_1_x_locator1);
  gfmult gfm_alpha369_2_x_locator2(10'b0101100101, locator2, alpha369_2_x_locator2);
  gfmult gfm_alpha369_3_x_locator3(10'b0111000100, locator3, alpha369_3_x_locator3);
  gfmult gfm_alpha370_0_x_locator0(10'b0000000001, locator0, alpha370_0_x_locator0);
  gfmult gfm_alpha370_1_x_locator1(10'b1000101000, locator1, alpha370_1_x_locator1);
  gfmult gfm_alpha370_2_x_locator2(10'b0101011011, locator2, alpha370_2_x_locator2);
  gfmult gfm_alpha370_3_x_locator3(10'b1000111100, locator3, alpha370_3_x_locator3);
  gfmult gfm_alpha371_0_x_locator0(10'b0000000001, locator0, alpha371_0_x_locator0);
  gfmult gfm_alpha371_1_x_locator1(10'b0100010100, locator1, alpha371_1_x_locator1);
  gfmult gfm_alpha371_2_x_locator2(10'b1101010000, locator2, alpha371_2_x_locator2);
  gfmult gfm_alpha371_3_x_locator3(10'b1001000011, locator3, alpha371_3_x_locator3);
  gfmult gfm_alpha372_0_x_locator0(10'b0000000001, locator0, alpha372_0_x_locator0);
  gfmult gfm_alpha372_1_x_locator1(10'b0010001010, locator1, alpha372_1_x_locator1);
  gfmult gfm_alpha372_2_x_locator2(10'b0011010100, locator2, alpha372_2_x_locator2);
  gfmult gfm_alpha372_3_x_locator3(10'b0111001011, locator3, alpha372_3_x_locator3);
  gfmult gfm_alpha373_0_x_locator0(10'b0000000001, locator0, alpha373_0_x_locator0);
  gfmult gfm_alpha373_1_x_locator1(10'b0001000101, locator1, alpha373_1_x_locator1);
  gfmult gfm_alpha373_2_x_locator2(10'b0000110101, locator2, alpha373_2_x_locator2);
  gfmult gfm_alpha373_3_x_locator3(10'b0110111010, locator3, alpha373_3_x_locator3);
  gfmult gfm_alpha374_0_x_locator0(10'b0000000001, locator0, alpha374_0_x_locator0);
  gfmult gfm_alpha374_1_x_locator1(10'b1000100110, locator1, alpha374_1_x_locator1);
  gfmult gfm_alpha374_2_x_locator2(10'b0100001111, locator2, alpha374_2_x_locator2);
  gfmult gfm_alpha374_3_x_locator3(10'b0100110101, locator3, alpha374_3_x_locator3);
  gfmult gfm_alpha375_0_x_locator0(10'b0000000001, locator0, alpha375_0_x_locator0);
  gfmult gfm_alpha375_1_x_locator1(10'b0100010011, locator1, alpha375_1_x_locator1);
  gfmult gfm_alpha375_2_x_locator2(10'b1101000101, locator2, alpha375_2_x_locator2);
  gfmult gfm_alpha375_3_x_locator3(10'b1010100011, locator3, alpha375_3_x_locator3);
  gfmult gfm_alpha376_0_x_locator0(10'b0000000001, locator0, alpha376_0_x_locator0);
  gfmult gfm_alpha376_1_x_locator1(10'b1010001101, locator1, alpha376_1_x_locator1);
  gfmult gfm_alpha376_2_x_locator2(10'b0111010011, locator2, alpha376_2_x_locator2);
  gfmult gfm_alpha376_3_x_locator3(10'b0111010111, locator3, alpha376_3_x_locator3);
  gfmult gfm_alpha377_0_x_locator0(10'b0000000001, locator0, alpha377_0_x_locator0);
  gfmult gfm_alpha377_1_x_locator1(10'b1101000010, locator1, alpha377_1_x_locator1);
  gfmult gfm_alpha377_2_x_locator2(10'b1101110010, locator2, alpha377_2_x_locator2);
  gfmult gfm_alpha377_3_x_locator3(10'b1110111101, locator3, alpha377_3_x_locator3);
  gfmult gfm_alpha378_0_x_locator0(10'b0000000001, locator0, alpha378_0_x_locator0);
  gfmult gfm_alpha378_1_x_locator1(10'b0110100001, locator1, alpha378_1_x_locator1);
  gfmult gfm_alpha378_2_x_locator2(10'b1011011000, locator2, alpha378_2_x_locator2);
  gfmult gfm_alpha378_3_x_locator3(10'b1011110010, locator3, alpha378_3_x_locator3);
  gfmult gfm_alpha379_0_x_locator0(10'b0000000001, locator0, alpha379_0_x_locator0);
  gfmult gfm_alpha379_1_x_locator1(10'b1011010100, locator1, alpha379_1_x_locator1);
  gfmult gfm_alpha379_2_x_locator2(10'b0010110110, locator2, alpha379_2_x_locator2);
  gfmult gfm_alpha379_3_x_locator3(10'b0101011100, locator3, alpha379_3_x_locator3);
  gfmult gfm_alpha380_0_x_locator0(10'b0000000001, locator0, alpha380_0_x_locator0);
  gfmult gfm_alpha380_1_x_locator1(10'b0101101010, locator1, alpha380_1_x_locator1);
  gfmult gfm_alpha380_2_x_locator2(10'b1000101001, locator2, alpha380_2_x_locator2);
  gfmult gfm_alpha380_3_x_locator3(10'b1000101111, locator3, alpha380_3_x_locator3);
  gfmult gfm_alpha381_0_x_locator0(10'b0000000001, locator0, alpha381_0_x_locator0);
  gfmult gfm_alpha381_1_x_locator1(10'b0010110101, locator1, alpha381_1_x_locator1);
  gfmult gfm_alpha381_2_x_locator2(10'b0110001000, locator2, alpha381_2_x_locator2);
  gfmult gfm_alpha381_3_x_locator3(10'b1111000010, locator3, alpha381_3_x_locator3);
  gfmult gfm_alpha382_0_x_locator0(10'b0000000001, locator0, alpha382_0_x_locator0);
  gfmult gfm_alpha382_1_x_locator1(10'b1001011110, locator1, alpha382_1_x_locator1);
  gfmult gfm_alpha382_2_x_locator2(10'b0001100010, locator2, alpha382_2_x_locator2);
  gfmult gfm_alpha382_3_x_locator3(10'b0101111010, locator3, alpha382_3_x_locator3);
  gfmult gfm_alpha383_0_x_locator0(10'b0000000001, locator0, alpha383_0_x_locator0);
  gfmult gfm_alpha383_1_x_locator1(10'b0100101111, locator1, alpha383_1_x_locator1);
  gfmult gfm_alpha383_2_x_locator2(10'b1000011100, locator2, alpha383_2_x_locator2);
  gfmult gfm_alpha383_3_x_locator3(10'b0100101101, locator3, alpha383_3_x_locator3);
  gfmult gfm_alpha384_0_x_locator0(10'b0000000001, locator0, alpha384_0_x_locator0);
  gfmult gfm_alpha384_1_x_locator1(10'b1010010011, locator1, alpha384_1_x_locator1);
  gfmult gfm_alpha384_2_x_locator2(10'b0010000111, locator2, alpha384_2_x_locator2);
  gfmult gfm_alpha384_3_x_locator3(10'b1010100000, locator3, alpha384_3_x_locator3);
  gfmult gfm_alpha385_0_x_locator0(10'b0000000001, locator0, alpha385_0_x_locator0);
  gfmult gfm_alpha385_1_x_locator1(10'b1101001101, locator1, alpha385_1_x_locator1);
  gfmult gfm_alpha385_2_x_locator2(10'b1100100111, locator2, alpha385_2_x_locator2);
  gfmult gfm_alpha385_3_x_locator3(10'b0001010100, locator3, alpha385_3_x_locator3);
  gfmult gfm_alpha386_0_x_locator0(10'b0000000001, locator0, alpha386_0_x_locator0);
  gfmult gfm_alpha386_1_x_locator1(10'b1110100010, locator1, alpha386_1_x_locator1);
  gfmult gfm_alpha386_2_x_locator2(10'b1111001111, locator2, alpha386_2_x_locator2);
  gfmult gfm_alpha386_3_x_locator3(10'b1000001110, locator3, alpha386_3_x_locator3);
  gfmult gfm_alpha387_0_x_locator0(10'b0000000001, locator0, alpha387_0_x_locator0);
  gfmult gfm_alpha387_1_x_locator1(10'b0111010001, locator1, alpha387_1_x_locator1);
  gfmult gfm_alpha387_2_x_locator2(10'b1111110101, locator2, alpha387_2_x_locator2);
  gfmult gfm_alpha387_3_x_locator3(10'b1101000111, locator3, alpha387_3_x_locator3);
  gfmult gfm_alpha388_0_x_locator0(10'b0000000001, locator0, alpha388_0_x_locator0);
  gfmult gfm_alpha388_1_x_locator1(10'b1011101100, locator1, alpha388_1_x_locator1);
  gfmult gfm_alpha388_2_x_locator2(10'b0111111111, locator2, alpha388_2_x_locator2);
  gfmult gfm_alpha388_3_x_locator3(10'b1111101111, locator3, alpha388_3_x_locator3);
  gfmult gfm_alpha389_0_x_locator0(10'b0000000001, locator0, alpha389_0_x_locator0);
  gfmult gfm_alpha389_1_x_locator1(10'b0101110110, locator1, alpha389_1_x_locator1);
  gfmult gfm_alpha389_2_x_locator2(10'b1101111001, locator2, alpha389_2_x_locator2);
  gfmult gfm_alpha389_3_x_locator3(10'b1111111010, locator3, alpha389_3_x_locator3);
  gfmult gfm_alpha390_0_x_locator0(10'b0000000001, locator0, alpha390_0_x_locator0);
  gfmult gfm_alpha390_1_x_locator1(10'b0010111011, locator1, alpha390_1_x_locator1);
  gfmult gfm_alpha390_2_x_locator2(10'b0111011100, locator2, alpha390_2_x_locator2);
  gfmult gfm_alpha390_3_x_locator3(10'b0101111101, locator3, alpha390_3_x_locator3);
  gfmult gfm_alpha391_0_x_locator0(10'b0000000001, locator0, alpha391_0_x_locator0);
  gfmult gfm_alpha391_1_x_locator1(10'b1001011001, locator1, alpha391_1_x_locator1);
  gfmult gfm_alpha391_2_x_locator2(10'b0001110111, locator2, alpha391_2_x_locator2);
  gfmult gfm_alpha391_3_x_locator3(10'b1010101010, locator3, alpha391_3_x_locator3);
  gfmult gfm_alpha392_0_x_locator0(10'b0000000001, locator0, alpha392_0_x_locator0);
  gfmult gfm_alpha392_1_x_locator1(10'b1100101000, locator1, alpha392_1_x_locator1);
  gfmult gfm_alpha392_2_x_locator2(10'b1100011011, locator2, alpha392_2_x_locator2);
  gfmult gfm_alpha392_3_x_locator3(10'b0101010111, locator3, alpha392_3_x_locator3);
  gfmult gfm_alpha393_0_x_locator0(10'b0000000001, locator0, alpha393_0_x_locator0);
  gfmult gfm_alpha393_1_x_locator1(10'b0110010100, locator1, alpha393_1_x_locator1);
  gfmult gfm_alpha393_2_x_locator2(10'b1111000000, locator2, alpha393_2_x_locator2);
  gfmult gfm_alpha393_3_x_locator3(10'b1110101101, locator3, alpha393_3_x_locator3);
  gfmult gfm_alpha394_0_x_locator0(10'b0000000001, locator0, alpha394_0_x_locator0);
  gfmult gfm_alpha394_1_x_locator1(10'b0011001010, locator1, alpha394_1_x_locator1);
  gfmult gfm_alpha394_2_x_locator2(10'b0011110000, locator2, alpha394_2_x_locator2);
  gfmult gfm_alpha394_3_x_locator3(10'b1011110000, locator3, alpha394_3_x_locator3);
  gfmult gfm_alpha395_0_x_locator0(10'b0000000001, locator0, alpha395_0_x_locator0);
  gfmult gfm_alpha395_1_x_locator1(10'b0001100101, locator1, alpha395_1_x_locator1);
  gfmult gfm_alpha395_2_x_locator2(10'b0000111100, locator2, alpha395_2_x_locator2);
  gfmult gfm_alpha395_3_x_locator3(10'b0001011110, locator3, alpha395_3_x_locator3);
  gfmult gfm_alpha396_0_x_locator0(10'b0000000001, locator0, alpha396_0_x_locator0);
  gfmult gfm_alpha396_1_x_locator1(10'b1000110110, locator1, alpha396_1_x_locator1);
  gfmult gfm_alpha396_2_x_locator2(10'b0000001111, locator2, alpha396_2_x_locator2);
  gfmult gfm_alpha396_3_x_locator3(10'b1100001101, locator3, alpha396_3_x_locator3);
  gfmult gfm_alpha397_0_x_locator0(10'b0000000001, locator0, alpha397_0_x_locator0);
  gfmult gfm_alpha397_1_x_locator1(10'b0100011011, locator1, alpha397_1_x_locator1);
  gfmult gfm_alpha397_2_x_locator2(10'b1100000101, locator2, alpha397_2_x_locator2);
  gfmult gfm_alpha397_3_x_locator3(10'b1011100100, locator3, alpha397_3_x_locator3);
  gfmult gfm_alpha398_0_x_locator0(10'b0000000001, locator0, alpha398_0_x_locator0);
  gfmult gfm_alpha398_1_x_locator1(10'b1010001001, locator1, alpha398_1_x_locator1);
  gfmult gfm_alpha398_2_x_locator2(10'b0111000011, locator2, alpha398_2_x_locator2);
  gfmult gfm_alpha398_3_x_locator3(10'b1001011000, locator3, alpha398_3_x_locator3);
  gfmult gfm_alpha399_0_x_locator0(10'b0000000001, locator0, alpha399_0_x_locator0);
  gfmult gfm_alpha399_1_x_locator1(10'b1101000000, locator1, alpha399_1_x_locator1);
  gfmult gfm_alpha399_2_x_locator2(10'b1101110110, locator2, alpha399_2_x_locator2);
  gfmult gfm_alpha399_3_x_locator3(10'b0001001011, locator3, alpha399_3_x_locator3);
  gfmult gfm_alpha400_0_x_locator0(10'b0000000001, locator0, alpha400_0_x_locator0);
  gfmult gfm_alpha400_1_x_locator1(10'b0110100000, locator1, alpha400_1_x_locator1);
  gfmult gfm_alpha400_2_x_locator2(10'b1011011001, locator2, alpha400_2_x_locator2);
  gfmult gfm_alpha400_3_x_locator3(10'b0110001010, locator3, alpha400_3_x_locator3);
  gfmult gfm_alpha401_0_x_locator0(10'b0000000001, locator0, alpha401_0_x_locator0);
  gfmult gfm_alpha401_1_x_locator1(10'b0011010000, locator1, alpha401_1_x_locator1);
  gfmult gfm_alpha401_2_x_locator2(10'b0110110100, locator2, alpha401_2_x_locator2);
  gfmult gfm_alpha401_3_x_locator3(10'b0100110011, locator3, alpha401_3_x_locator3);
  gfmult gfm_alpha402_0_x_locator0(10'b0000000001, locator0, alpha402_0_x_locator0);
  gfmult gfm_alpha402_1_x_locator1(10'b0001101000, locator1, alpha402_1_x_locator1);
  gfmult gfm_alpha402_2_x_locator2(10'b0001101101, locator2, alpha402_2_x_locator2);
  gfmult gfm_alpha402_3_x_locator3(10'b0110100101, locator3, alpha402_3_x_locator3);
  gfmult gfm_alpha403_0_x_locator0(10'b0000000001, locator0, alpha403_0_x_locator0);
  gfmult gfm_alpha403_1_x_locator1(10'b0000110100, locator1, alpha403_1_x_locator1);
  gfmult gfm_alpha403_2_x_locator2(10'b0100011001, locator2, alpha403_2_x_locator2);
  gfmult gfm_alpha403_3_x_locator3(10'b1010110001, locator3, alpha403_3_x_locator3);
  gfmult gfm_alpha404_0_x_locator0(10'b0000000001, locator0, alpha404_0_x_locator0);
  gfmult gfm_alpha404_1_x_locator1(10'b0000011010, locator1, alpha404_1_x_locator1);
  gfmult gfm_alpha404_2_x_locator2(10'b0101000100, locator2, alpha404_2_x_locator2);
  gfmult gfm_alpha404_3_x_locator3(10'b0011010111, locator3, alpha404_3_x_locator3);
  gfmult gfm_alpha405_0_x_locator0(10'b0000000001, locator0, alpha405_0_x_locator0);
  gfmult gfm_alpha405_1_x_locator1(10'b0000001101, locator1, alpha405_1_x_locator1);
  gfmult gfm_alpha405_2_x_locator2(10'b0001010001, locator2, alpha405_2_x_locator2);
  gfmult gfm_alpha405_3_x_locator3(10'b1110011101, locator3, alpha405_3_x_locator3);
  gfmult gfm_alpha406_0_x_locator0(10'b0000000001, locator0, alpha406_0_x_locator0);
  gfmult gfm_alpha406_1_x_locator1(10'b1000000010, locator1, alpha406_1_x_locator1);
  gfmult gfm_alpha406_2_x_locator2(10'b0100010110, locator2, alpha406_2_x_locator2);
  gfmult gfm_alpha406_3_x_locator3(10'b1011110110, locator3, alpha406_3_x_locator3);
  gfmult gfm_alpha407_0_x_locator0(10'b0000000001, locator0, alpha407_0_x_locator0);
  gfmult gfm_alpha407_1_x_locator1(10'b0100000001, locator1, alpha407_1_x_locator1);
  gfmult gfm_alpha407_2_x_locator2(10'b1001000001, locator2, alpha407_2_x_locator2);
  gfmult gfm_alpha407_3_x_locator3(10'b1101011000, locator3, alpha407_3_x_locator3);
  gfmult gfm_alpha408_0_x_locator0(10'b0000000001, locator0, alpha408_0_x_locator0);
  gfmult gfm_alpha408_1_x_locator1(10'b1010000100, locator1, alpha408_1_x_locator1);
  gfmult gfm_alpha408_2_x_locator2(10'b0110010010, locator2, alpha408_2_x_locator2);
  gfmult gfm_alpha408_3_x_locator3(10'b0001101011, locator3, alpha408_3_x_locator3);
  gfmult gfm_alpha409_0_x_locator0(10'b0000000001, locator0, alpha409_0_x_locator0);
  gfmult gfm_alpha409_1_x_locator1(10'b0101000010, locator1, alpha409_1_x_locator1);
  gfmult gfm_alpha409_2_x_locator2(10'b1001100000, locator2, alpha409_2_x_locator2);
  gfmult gfm_alpha409_3_x_locator3(10'b0110001110, locator3, alpha409_3_x_locator3);
  gfmult gfm_alpha410_0_x_locator0(10'b0000000001, locator0, alpha410_0_x_locator0);
  gfmult gfm_alpha410_1_x_locator1(10'b0010100001, locator1, alpha410_1_x_locator1);
  gfmult gfm_alpha410_2_x_locator2(10'b0010011000, locator2, alpha410_2_x_locator2);
  gfmult gfm_alpha410_3_x_locator3(10'b1100110111, locator3, alpha410_3_x_locator3);
  gfmult gfm_alpha411_0_x_locator0(10'b0000000001, locator0, alpha411_0_x_locator0);
  gfmult gfm_alpha411_1_x_locator1(10'b1001010100, locator1, alpha411_1_x_locator1);
  gfmult gfm_alpha411_2_x_locator2(10'b0000100110, locator2, alpha411_2_x_locator2);
  gfmult gfm_alpha411_3_x_locator3(10'b1111100001, locator3, alpha411_3_x_locator3);
  gfmult gfm_alpha412_0_x_locator0(10'b0000000001, locator0, alpha412_0_x_locator0);
  gfmult gfm_alpha412_1_x_locator1(10'b0100101010, locator1, alpha412_1_x_locator1);
  gfmult gfm_alpha412_2_x_locator2(10'b1000001101, locator2, alpha412_2_x_locator2);
  gfmult gfm_alpha412_3_x_locator3(10'b0011111101, locator3, alpha412_3_x_locator3);
  gfmult gfm_alpha413_0_x_locator0(10'b0000000001, locator0, alpha413_0_x_locator0);
  gfmult gfm_alpha413_1_x_locator1(10'b0010010101, locator1, alpha413_1_x_locator1);
  gfmult gfm_alpha413_2_x_locator2(10'b0110000001, locator2, alpha413_2_x_locator2);
  gfmult gfm_alpha413_3_x_locator3(10'b1010011010, locator3, alpha413_3_x_locator3);
  gfmult gfm_alpha414_0_x_locator0(10'b0000000001, locator0, alpha414_0_x_locator0);
  gfmult gfm_alpha414_1_x_locator1(10'b1001001110, locator1, alpha414_1_x_locator1);
  gfmult gfm_alpha414_2_x_locator2(10'b0101100010, locator2, alpha414_2_x_locator2);
  gfmult gfm_alpha414_3_x_locator3(10'b0101010001, locator3, alpha414_3_x_locator3);
  gfmult gfm_alpha415_0_x_locator0(10'b0000000001, locator0, alpha415_0_x_locator0);
  gfmult gfm_alpha415_1_x_locator1(10'b0100100111, locator1, alpha415_1_x_locator1);
  gfmult gfm_alpha415_2_x_locator2(10'b1001011100, locator2, alpha415_2_x_locator2);
  gfmult gfm_alpha415_3_x_locator3(10'b0010101011, locator3, alpha415_3_x_locator3);
  gfmult gfm_alpha416_0_x_locator0(10'b0000000001, locator0, alpha416_0_x_locator0);
  gfmult gfm_alpha416_1_x_locator1(10'b1010010111, locator1, alpha416_1_x_locator1);
  gfmult gfm_alpha416_2_x_locator2(10'b0010010111, locator2, alpha416_2_x_locator2);
  gfmult gfm_alpha416_3_x_locator3(10'b0110010110, locator3, alpha416_3_x_locator3);
  gfmult gfm_alpha417_0_x_locator0(10'b0000000001, locator0, alpha417_0_x_locator0);
  gfmult gfm_alpha417_1_x_locator1(10'b1101001111, locator1, alpha417_1_x_locator1);
  gfmult gfm_alpha417_2_x_locator2(10'b1100100011, locator2, alpha417_2_x_locator2);
  gfmult gfm_alpha417_3_x_locator3(10'b1100110100, locator3, alpha417_3_x_locator3);
  gfmult gfm_alpha418_0_x_locator0(10'b0000000001, locator0, alpha418_0_x_locator0);
  gfmult gfm_alpha418_1_x_locator1(10'b1110100011, locator1, alpha418_1_x_locator1);
  gfmult gfm_alpha418_2_x_locator2(10'b1111001110, locator2, alpha418_2_x_locator2);
  gfmult gfm_alpha418_3_x_locator3(10'b1001100010, locator3, alpha418_3_x_locator3);
  gfmult gfm_alpha419_0_x_locator0(10'b0000000001, locator0, alpha419_0_x_locator0);
  gfmult gfm_alpha419_1_x_locator1(10'b1111010101, locator1, alpha419_1_x_locator1);
  gfmult gfm_alpha419_2_x_locator2(10'b1011110111, locator2, alpha419_2_x_locator2);
  gfmult gfm_alpha419_3_x_locator3(10'b0101001110, locator3, alpha419_3_x_locator3);
  gfmult gfm_alpha420_0_x_locator0(10'b0000000001, locator0, alpha420_0_x_locator0);
  gfmult gfm_alpha420_1_x_locator1(10'b1111101110, locator1, alpha420_1_x_locator1);
  gfmult gfm_alpha420_2_x_locator2(10'b1110111011, locator2, alpha420_2_x_locator2);
  gfmult gfm_alpha420_3_x_locator3(10'b1100101111, locator3, alpha420_3_x_locator3);
  gfmult gfm_alpha421_0_x_locator0(10'b0000000001, locator0, alpha421_0_x_locator0);
  gfmult gfm_alpha421_1_x_locator1(10'b0111110111, locator1, alpha421_1_x_locator1);
  gfmult gfm_alpha421_2_x_locator2(10'b1111101000, locator2, alpha421_2_x_locator2);
  gfmult gfm_alpha421_3_x_locator3(10'b1111100010, locator3, alpha421_3_x_locator3);
  gfmult gfm_alpha422_0_x_locator0(10'b0000000001, locator0, alpha422_0_x_locator0);
  gfmult gfm_alpha422_1_x_locator1(10'b1011111111, locator1, alpha422_1_x_locator1);
  gfmult gfm_alpha422_2_x_locator2(10'b0011111010, locator2, alpha422_2_x_locator2);
  gfmult gfm_alpha422_3_x_locator3(10'b0101111110, locator3, alpha422_3_x_locator3);
  gfmult gfm_alpha423_0_x_locator0(10'b0000000001, locator0, alpha423_0_x_locator0);
  gfmult gfm_alpha423_1_x_locator1(10'b1101111011, locator1, alpha423_1_x_locator1);
  gfmult gfm_alpha423_2_x_locator2(10'b1000111010, locator2, alpha423_2_x_locator2);
  gfmult gfm_alpha423_3_x_locator3(10'b1100101001, locator3, alpha423_3_x_locator3);
  gfmult gfm_alpha424_0_x_locator0(10'b0000000001, locator0, alpha424_0_x_locator0);
  gfmult gfm_alpha424_1_x_locator1(10'b1110111001, locator1, alpha424_1_x_locator1);
  gfmult gfm_alpha424_2_x_locator2(10'b1010001010, locator2, alpha424_2_x_locator2);
  gfmult gfm_alpha424_3_x_locator3(10'b0011100100, locator3, alpha424_3_x_locator3);
  gfmult gfm_alpha425_0_x_locator0(10'b0000000001, locator0, alpha425_0_x_locator0);
  gfmult gfm_alpha425_1_x_locator1(10'b1111011000, locator1, alpha425_1_x_locator1);
  gfmult gfm_alpha425_2_x_locator2(10'b1010100110, locator2, alpha425_2_x_locator2);
  gfmult gfm_alpha425_3_x_locator3(10'b1000011000, locator3, alpha425_3_x_locator3);
  gfmult gfm_alpha426_0_x_locator0(10'b0000000001, locator0, alpha426_0_x_locator0);
  gfmult gfm_alpha426_1_x_locator1(10'b0111101100, locator1, alpha426_1_x_locator1);
  gfmult gfm_alpha426_2_x_locator2(10'b1010101101, locator2, alpha426_2_x_locator2);
  gfmult gfm_alpha426_3_x_locator3(10'b0001000011, locator3, alpha426_3_x_locator3);
  gfmult gfm_alpha427_0_x_locator0(10'b0000000001, locator0, alpha427_0_x_locator0);
  gfmult gfm_alpha427_1_x_locator1(10'b0011110110, locator1, alpha427_1_x_locator1);
  gfmult gfm_alpha427_2_x_locator2(10'b0110101001, locator2, alpha427_2_x_locator2);
  gfmult gfm_alpha427_3_x_locator3(10'b0110001011, locator3, alpha427_3_x_locator3);
  gfmult gfm_alpha428_0_x_locator0(10'b0000000001, locator0, alpha428_0_x_locator0);
  gfmult gfm_alpha428_1_x_locator1(10'b0001111011, locator1, alpha428_1_x_locator1);
  gfmult gfm_alpha428_2_x_locator2(10'b0101101000, locator2, alpha428_2_x_locator2);
  gfmult gfm_alpha428_3_x_locator3(10'b0110110010, locator3, alpha428_3_x_locator3);
  gfmult gfm_alpha429_0_x_locator0(10'b0000000001, locator0, alpha429_0_x_locator0);
  gfmult gfm_alpha429_1_x_locator1(10'b1000111001, locator1, alpha429_1_x_locator1);
  gfmult gfm_alpha429_2_x_locator2(10'b0001011010, locator2, alpha429_2_x_locator2);
  gfmult gfm_alpha429_3_x_locator3(10'b0100110100, locator3, alpha429_3_x_locator3);
  gfmult gfm_alpha430_0_x_locator0(10'b0000000001, locator0, alpha430_0_x_locator0);
  gfmult gfm_alpha430_1_x_locator1(10'b1100011000, locator1, alpha430_1_x_locator1);
  gfmult gfm_alpha430_2_x_locator2(10'b1000010010, locator2, alpha430_2_x_locator2);
  gfmult gfm_alpha430_3_x_locator3(10'b1000100010, locator3, alpha430_3_x_locator3);
  gfmult gfm_alpha431_0_x_locator0(10'b0000000001, locator0, alpha431_0_x_locator0);
  gfmult gfm_alpha431_1_x_locator1(10'b0110001100, locator1, alpha431_1_x_locator1);
  gfmult gfm_alpha431_2_x_locator2(10'b1010000000, locator2, alpha431_2_x_locator2);
  gfmult gfm_alpha431_3_x_locator3(10'b0101000110, locator3, alpha431_3_x_locator3);
  gfmult gfm_alpha432_0_x_locator0(10'b0000000001, locator0, alpha432_0_x_locator0);
  gfmult gfm_alpha432_1_x_locator1(10'b0011000110, locator1, alpha432_1_x_locator1);
  gfmult gfm_alpha432_2_x_locator2(10'b0010100000, locator2, alpha432_2_x_locator2);
  gfmult gfm_alpha432_3_x_locator3(10'b1100101110, locator3, alpha432_3_x_locator3);
  gfmult gfm_alpha433_0_x_locator0(10'b0000000001, locator0, alpha433_0_x_locator0);
  gfmult gfm_alpha433_1_x_locator1(10'b0001100011, locator1, alpha433_1_x_locator1);
  gfmult gfm_alpha433_2_x_locator2(10'b0000101000, locator2, alpha433_2_x_locator2);
  gfmult gfm_alpha433_3_x_locator3(10'b1101100011, locator3, alpha433_3_x_locator3);
  gfmult gfm_alpha434_0_x_locator0(10'b0000000001, locator0, alpha434_0_x_locator0);
  gfmult gfm_alpha434_1_x_locator1(10'b1000110101, locator1, alpha434_1_x_locator1);
  gfmult gfm_alpha434_2_x_locator2(10'b0000001010, locator2, alpha434_2_x_locator2);
  gfmult gfm_alpha434_3_x_locator3(10'b0111101111, locator3, alpha434_3_x_locator3);
  gfmult gfm_alpha435_0_x_locator0(10'b0000000001, locator0, alpha435_0_x_locator0);
  gfmult gfm_alpha435_1_x_locator1(10'b1100011110, locator1, alpha435_1_x_locator1);
  gfmult gfm_alpha435_2_x_locator2(10'b1000000110, locator2, alpha435_2_x_locator2);
  gfmult gfm_alpha435_3_x_locator3(10'b1110111010, locator3, alpha435_3_x_locator3);
  gfmult gfm_alpha436_0_x_locator0(10'b0000000001, locator0, alpha436_0_x_locator0);
  gfmult gfm_alpha436_1_x_locator1(10'b0110001111, locator1, alpha436_1_x_locator1);
  gfmult gfm_alpha436_2_x_locator2(10'b1010000101, locator2, alpha436_2_x_locator2);
  gfmult gfm_alpha436_3_x_locator3(10'b0101110101, locator3, alpha436_3_x_locator3);
  gfmult gfm_alpha437_0_x_locator0(10'b0000000001, locator0, alpha437_0_x_locator0);
  gfmult gfm_alpha437_1_x_locator1(10'b1011000011, locator1, alpha437_1_x_locator1);
  gfmult gfm_alpha437_2_x_locator2(10'b0110100011, locator2, alpha437_2_x_locator2);
  gfmult gfm_alpha437_3_x_locator3(10'b1010101011, locator3, alpha437_3_x_locator3);
  gfmult gfm_alpha438_0_x_locator0(10'b0000000001, locator0, alpha438_0_x_locator0);
  gfmult gfm_alpha438_1_x_locator1(10'b1101100101, locator1, alpha438_1_x_locator1);
  gfmult gfm_alpha438_2_x_locator2(10'b1101101110, locator2, alpha438_2_x_locator2);
  gfmult gfm_alpha438_3_x_locator3(10'b0111010110, locator3, alpha438_3_x_locator3);
  gfmult gfm_alpha439_0_x_locator0(10'b0000000001, locator0, alpha439_0_x_locator0);
  gfmult gfm_alpha439_1_x_locator1(10'b1110110110, locator1, alpha439_1_x_locator1);
  gfmult gfm_alpha439_2_x_locator2(10'b1011011111, locator2, alpha439_2_x_locator2);
  gfmult gfm_alpha439_3_x_locator3(10'b1100111100, locator3, alpha439_3_x_locator3);
  gfmult gfm_alpha440_0_x_locator0(10'b0000000001, locator0, alpha440_0_x_locator0);
  gfmult gfm_alpha440_1_x_locator1(10'b0111011011, locator1, alpha440_1_x_locator1);
  gfmult gfm_alpha440_2_x_locator2(10'b1110110001, locator2, alpha440_2_x_locator2);
  gfmult gfm_alpha440_3_x_locator3(10'b1001100011, locator3, alpha440_3_x_locator3);
  gfmult gfm_alpha441_0_x_locator0(10'b0000000001, locator0, alpha441_0_x_locator0);
  gfmult gfm_alpha441_1_x_locator1(10'b1011101001, locator1, alpha441_1_x_locator1);
  gfmult gfm_alpha441_2_x_locator2(10'b0111101110, locator2, alpha441_2_x_locator2);
  gfmult gfm_alpha441_3_x_locator3(10'b0111001111, locator3, alpha441_3_x_locator3);
  gfmult gfm_alpha442_0_x_locator0(10'b0000000001, locator0, alpha442_0_x_locator0);
  gfmult gfm_alpha442_1_x_locator1(10'b1101110000, locator1, alpha442_1_x_locator1);
  gfmult gfm_alpha442_2_x_locator2(10'b1001111111, locator2, alpha442_2_x_locator2);
  gfmult gfm_alpha442_3_x_locator3(10'b1110111110, locator3, alpha442_3_x_locator3);
  gfmult gfm_alpha443_0_x_locator0(10'b0000000001, locator0, alpha443_0_x_locator0);
  gfmult gfm_alpha443_1_x_locator1(10'b0110111000, locator1, alpha443_1_x_locator1);
  gfmult gfm_alpha443_2_x_locator2(10'b1110011001, locator2, alpha443_2_x_locator2);
  gfmult gfm_alpha443_3_x_locator3(10'b1101110001, locator3, alpha443_3_x_locator3);
  gfmult gfm_alpha444_0_x_locator0(10'b0000000001, locator0, alpha444_0_x_locator0);
  gfmult gfm_alpha444_1_x_locator1(10'b0011011100, locator1, alpha444_1_x_locator1);
  gfmult gfm_alpha444_2_x_locator2(10'b0111100100, locator2, alpha444_2_x_locator2);
  gfmult gfm_alpha444_3_x_locator3(10'b0011101111, locator3, alpha444_3_x_locator3);
  gfmult gfm_alpha445_0_x_locator0(10'b0000000001, locator0, alpha445_0_x_locator0);
  gfmult gfm_alpha445_1_x_locator1(10'b0001101110, locator1, alpha445_1_x_locator1);
  gfmult gfm_alpha445_2_x_locator2(10'b0001111001, locator2, alpha445_2_x_locator2);
  gfmult gfm_alpha445_3_x_locator3(10'b1110011010, locator3, alpha445_3_x_locator3);
  gfmult gfm_alpha446_0_x_locator0(10'b0000000001, locator0, alpha446_0_x_locator0);
  gfmult gfm_alpha446_1_x_locator1(10'b0000110111, locator1, alpha446_1_x_locator1);
  gfmult gfm_alpha446_2_x_locator2(10'b0100011100, locator2, alpha446_2_x_locator2);
  gfmult gfm_alpha446_3_x_locator3(10'b0101110001, locator3, alpha446_3_x_locator3);
  gfmult gfm_alpha447_0_x_locator0(10'b0000000001, locator0, alpha447_0_x_locator0);
  gfmult gfm_alpha447_1_x_locator1(10'b1000011111, locator1, alpha447_1_x_locator1);
  gfmult gfm_alpha447_2_x_locator2(10'b0001000111, locator2, alpha447_2_x_locator2);
  gfmult gfm_alpha447_3_x_locator3(10'b0010101111, locator3, alpha447_3_x_locator3);
  gfmult gfm_alpha448_0_x_locator0(10'b0000000001, locator0, alpha448_0_x_locator0);
  gfmult gfm_alpha448_1_x_locator1(10'b1100001011, locator1, alpha448_1_x_locator1);
  gfmult gfm_alpha448_2_x_locator2(10'b1100010111, locator2, alpha448_2_x_locator2);
  gfmult gfm_alpha448_3_x_locator3(10'b1110010010, locator3, alpha448_3_x_locator3);
  gfmult gfm_alpha449_0_x_locator0(10'b0000000001, locator0, alpha449_0_x_locator0);
  gfmult gfm_alpha449_1_x_locator1(10'b1110000001, locator1, alpha449_1_x_locator1);
  gfmult gfm_alpha449_2_x_locator2(10'b1111000011, locator2, alpha449_2_x_locator2);
  gfmult gfm_alpha449_3_x_locator3(10'b0101110000, locator3, alpha449_3_x_locator3);
  gfmult gfm_alpha450_0_x_locator0(10'b0000000001, locator0, alpha450_0_x_locator0);
  gfmult gfm_alpha450_1_x_locator1(10'b1111000100, locator1, alpha450_1_x_locator1);
  gfmult gfm_alpha450_2_x_locator2(10'b1111110110, locator2, alpha450_2_x_locator2);
  gfmult gfm_alpha450_3_x_locator3(10'b0000101110, locator3, alpha450_3_x_locator3);
  gfmult gfm_alpha451_0_x_locator0(10'b0000000001, locator0, alpha451_0_x_locator0);
  gfmult gfm_alpha451_1_x_locator1(10'b0111100010, locator1, alpha451_1_x_locator1);
  gfmult gfm_alpha451_2_x_locator2(10'b1011111001, locator2, alpha451_2_x_locator2);
  gfmult gfm_alpha451_3_x_locator3(10'b1100000011, locator3, alpha451_3_x_locator3);
  gfmult gfm_alpha452_0_x_locator0(10'b0000000001, locator0, alpha452_0_x_locator0);
  gfmult gfm_alpha452_1_x_locator1(10'b0011110001, locator1, alpha452_1_x_locator1);
  gfmult gfm_alpha452_2_x_locator2(10'b0110111100, locator2, alpha452_2_x_locator2);
  gfmult gfm_alpha452_3_x_locator3(10'b0111100011, locator3, alpha452_3_x_locator3);
  gfmult gfm_alpha453_0_x_locator0(10'b0000000001, locator0, alpha453_0_x_locator0);
  gfmult gfm_alpha453_1_x_locator1(10'b1001111100, locator1, alpha453_1_x_locator1);
  gfmult gfm_alpha453_2_x_locator2(10'b0001101111, locator2, alpha453_2_x_locator2);
  gfmult gfm_alpha453_3_x_locator3(10'b0110111111, locator3, alpha453_3_x_locator3);
  gfmult gfm_alpha454_0_x_locator0(10'b0000000001, locator0, alpha454_0_x_locator0);
  gfmult gfm_alpha454_1_x_locator1(10'b0100111110, locator1, alpha454_1_x_locator1);
  gfmult gfm_alpha454_2_x_locator2(10'b1100011101, locator2, alpha454_2_x_locator2);
  gfmult gfm_alpha454_3_x_locator3(10'b1110110000, locator3, alpha454_3_x_locator3);
  gfmult gfm_alpha455_0_x_locator0(10'b0000000001, locator0, alpha455_0_x_locator0);
  gfmult gfm_alpha455_1_x_locator1(10'b0010011111, locator1, alpha455_1_x_locator1);
  gfmult gfm_alpha455_2_x_locator2(10'b0111000101, locator2, alpha455_2_x_locator2);
  gfmult gfm_alpha455_3_x_locator3(10'b0001110110, locator3, alpha455_3_x_locator3);
  gfmult gfm_alpha456_0_x_locator0(10'b0000000001, locator0, alpha456_0_x_locator0);
  gfmult gfm_alpha456_1_x_locator1(10'b1001001011, locator1, alpha456_1_x_locator1);
  gfmult gfm_alpha456_2_x_locator2(10'b0101110011, locator2, alpha456_2_x_locator2);
  gfmult gfm_alpha456_3_x_locator3(10'b1100001000, locator3, alpha456_3_x_locator3);
  gfmult gfm_alpha457_0_x_locator0(10'b0000000001, locator0, alpha457_0_x_locator0);
  gfmult gfm_alpha457_1_x_locator1(10'b1100100001, locator1, alpha457_1_x_locator1);
  gfmult gfm_alpha457_2_x_locator2(10'b1101011010, locator2, alpha457_2_x_locator2);
  gfmult gfm_alpha457_3_x_locator3(10'b0001100001, locator3, alpha457_3_x_locator3);
  gfmult gfm_alpha458_0_x_locator0(10'b0000000001, locator0, alpha458_0_x_locator0);
  gfmult gfm_alpha458_1_x_locator1(10'b1110010100, locator1, alpha458_1_x_locator1);
  gfmult gfm_alpha458_2_x_locator2(10'b1011010010, locator2, alpha458_2_x_locator2);
  gfmult gfm_alpha458_3_x_locator3(10'b0010001101, locator3, alpha458_3_x_locator3);
  gfmult gfm_alpha459_0_x_locator0(10'b0000000001, locator0, alpha459_0_x_locator0);
  gfmult gfm_alpha459_1_x_locator1(10'b0111001010, locator1, alpha459_1_x_locator1);
  gfmult gfm_alpha459_2_x_locator2(10'b1010110000, locator2, alpha459_2_x_locator2);
  gfmult gfm_alpha459_3_x_locator3(10'b1010010100, locator3, alpha459_3_x_locator3);
  gfmult gfm_alpha460_0_x_locator0(10'b0000000001, locator0, alpha460_0_x_locator0);
  gfmult gfm_alpha460_1_x_locator1(10'b0011100101, locator1, alpha460_1_x_locator1);
  gfmult gfm_alpha460_2_x_locator2(10'b0010101100, locator2, alpha460_2_x_locator2);
  gfmult gfm_alpha460_3_x_locator3(10'b1001010110, locator3, alpha460_3_x_locator3);
  gfmult gfm_alpha461_0_x_locator0(10'b0000000001, locator0, alpha461_0_x_locator0);
  gfmult gfm_alpha461_1_x_locator1(10'b1001110110, locator1, alpha461_1_x_locator1);
  gfmult gfm_alpha461_2_x_locator2(10'b0000101011, locator2, alpha461_2_x_locator2);
  gfmult gfm_alpha461_3_x_locator3(10'b1101001100, locator3, alpha461_3_x_locator3);
  gfmult gfm_alpha462_0_x_locator0(10'b0000000001, locator0, alpha462_0_x_locator0);
  gfmult gfm_alpha462_1_x_locator1(10'b0100111011, locator1, alpha462_1_x_locator1);
  gfmult gfm_alpha462_2_x_locator2(10'b1100001100, locator2, alpha462_2_x_locator2);
  gfmult gfm_alpha462_3_x_locator3(10'b1001101101, locator3, alpha462_3_x_locator3);
  gfmult gfm_alpha463_0_x_locator0(10'b0000000001, locator0, alpha463_0_x_locator0);
  gfmult gfm_alpha463_1_x_locator1(10'b1010011001, locator1, alpha463_1_x_locator1);
  gfmult gfm_alpha463_2_x_locator2(10'b0011000011, locator2, alpha463_2_x_locator2);
  gfmult gfm_alpha463_3_x_locator3(10'b1011001000, locator3, alpha463_3_x_locator3);
  gfmult gfm_alpha464_0_x_locator0(10'b0000000001, locator0, alpha464_0_x_locator0);
  gfmult gfm_alpha464_1_x_locator1(10'b1101001000, locator1, alpha464_1_x_locator1);
  gfmult gfm_alpha464_2_x_locator2(10'b1100110110, locator2, alpha464_2_x_locator2);
  gfmult gfm_alpha464_3_x_locator3(10'b0001011001, locator3, alpha464_3_x_locator3);
  gfmult gfm_alpha465_0_x_locator0(10'b0000000001, locator0, alpha465_0_x_locator0);
  gfmult gfm_alpha465_1_x_locator1(10'b0110100100, locator1, alpha465_1_x_locator1);
  gfmult gfm_alpha465_2_x_locator2(10'b1011001001, locator2, alpha465_2_x_locator2);
  gfmult gfm_alpha465_3_x_locator3(10'b0010001010, locator3, alpha465_3_x_locator3);
  gfmult gfm_alpha466_0_x_locator0(10'b0000000001, locator0, alpha466_0_x_locator0);
  gfmult gfm_alpha466_1_x_locator1(10'b0011010010, locator1, alpha466_1_x_locator1);
  gfmult gfm_alpha466_2_x_locator2(10'b0110110000, locator2, alpha466_2_x_locator2);
  gfmult gfm_alpha466_3_x_locator3(10'b0100010011, locator3, alpha466_3_x_locator3);
  gfmult gfm_alpha467_0_x_locator0(10'b0000000001, locator0, alpha467_0_x_locator0);
  gfmult gfm_alpha467_1_x_locator1(10'b0001101001, locator1, alpha467_1_x_locator1);
  gfmult gfm_alpha467_2_x_locator2(10'b0001101100, locator2, alpha467_2_x_locator2);
  gfmult gfm_alpha467_3_x_locator3(10'b0110100001, locator3, alpha467_3_x_locator3);
  gfmult gfm_alpha468_0_x_locator0(10'b0000000001, locator0, alpha468_0_x_locator0);
  gfmult gfm_alpha468_1_x_locator1(10'b1000110000, locator1, alpha468_1_x_locator1);
  gfmult gfm_alpha468_2_x_locator2(10'b0000011011, locator2, alpha468_2_x_locator2);
  gfmult gfm_alpha468_3_x_locator3(10'b0010110101, locator3, alpha468_3_x_locator3);
  gfmult gfm_alpha469_0_x_locator0(10'b0000000001, locator0, alpha469_0_x_locator0);
  gfmult gfm_alpha469_1_x_locator1(10'b0100011000, locator1, alpha469_1_x_locator1);
  gfmult gfm_alpha469_2_x_locator2(10'b1100000000, locator2, alpha469_2_x_locator2);
  gfmult gfm_alpha469_3_x_locator3(10'b1010010011, locator3, alpha469_3_x_locator3);
  gfmult gfm_alpha470_0_x_locator0(10'b0000000001, locator0, alpha470_0_x_locator0);
  gfmult gfm_alpha470_1_x_locator1(10'b0010001100, locator1, alpha470_1_x_locator1);
  gfmult gfm_alpha470_2_x_locator2(10'b0011000000, locator2, alpha470_2_x_locator2);
  gfmult gfm_alpha470_3_x_locator3(10'b0111010001, locator3, alpha470_3_x_locator3);
  gfmult gfm_alpha471_0_x_locator0(10'b0000000001, locator0, alpha471_0_x_locator0);
  gfmult gfm_alpha471_1_x_locator1(10'b0001000110, locator1, alpha471_1_x_locator1);
  gfmult gfm_alpha471_2_x_locator2(10'b0000110000, locator2, alpha471_2_x_locator2);
  gfmult gfm_alpha471_3_x_locator3(10'b0010111011, locator3, alpha471_3_x_locator3);
  gfmult gfm_alpha472_0_x_locator0(10'b0000000001, locator0, alpha472_0_x_locator0);
  gfmult gfm_alpha472_1_x_locator1(10'b0000100011, locator1, alpha472_1_x_locator1);
  gfmult gfm_alpha472_2_x_locator2(10'b0000001100, locator2, alpha472_2_x_locator2);
  gfmult gfm_alpha472_3_x_locator3(10'b0110010100, locator3, alpha472_3_x_locator3);
  gfmult gfm_alpha473_0_x_locator0(10'b0000000001, locator0, alpha473_0_x_locator0);
  gfmult gfm_alpha473_1_x_locator1(10'b1000010101, locator1, alpha473_1_x_locator1);
  gfmult gfm_alpha473_2_x_locator2(10'b0000000011, locator2, alpha473_2_x_locator2);
  gfmult gfm_alpha473_3_x_locator3(10'b1000110110, locator3, alpha473_3_x_locator3);
  gfmult gfm_alpha474_0_x_locator0(10'b0000000001, locator0, alpha474_0_x_locator0);
  gfmult gfm_alpha474_1_x_locator1(10'b1100001110, locator1, alpha474_1_x_locator1);
  gfmult gfm_alpha474_2_x_locator2(10'b1100000110, locator2, alpha474_2_x_locator2);
  gfmult gfm_alpha474_3_x_locator3(10'b1101000000, locator3, alpha474_3_x_locator3);
  gfmult gfm_alpha475_0_x_locator0(10'b0000000001, locator0, alpha475_0_x_locator0);
  gfmult gfm_alpha475_1_x_locator1(10'b0110000111, locator1, alpha475_1_x_locator1);
  gfmult gfm_alpha475_2_x_locator2(10'b1011000101, locator2, alpha475_2_x_locator2);
  gfmult gfm_alpha475_3_x_locator3(10'b0001101000, locator3, alpha475_3_x_locator3);
  gfmult gfm_alpha476_0_x_locator0(10'b0000000001, locator0, alpha476_0_x_locator0);
  gfmult gfm_alpha476_1_x_locator1(10'b1011000111, locator1, alpha476_1_x_locator1);
  gfmult gfm_alpha476_2_x_locator2(10'b0110110011, locator2, alpha476_2_x_locator2);
  gfmult gfm_alpha476_3_x_locator3(10'b0000001101, locator3, alpha476_3_x_locator3);
  gfmult gfm_alpha477_0_x_locator0(10'b0000000001, locator0, alpha477_0_x_locator0);
  gfmult gfm_alpha477_1_x_locator1(10'b1101100111, locator1, alpha477_1_x_locator1);
  gfmult gfm_alpha477_2_x_locator2(10'b1101101010, locator2, alpha477_2_x_locator2);
  gfmult gfm_alpha477_3_x_locator3(10'b1010000100, locator3, alpha477_3_x_locator3);
  gfmult gfm_alpha478_0_x_locator0(10'b0000000001, locator0, alpha478_0_x_locator0);
  gfmult gfm_alpha478_1_x_locator1(10'b1110110111, locator1, alpha478_1_x_locator1);
  gfmult gfm_alpha478_2_x_locator2(10'b1011011110, locator2, alpha478_2_x_locator2);
  gfmult gfm_alpha478_3_x_locator3(10'b1001010100, locator3, alpha478_3_x_locator3);
  gfmult gfm_alpha479_0_x_locator0(10'b0000000001, locator0, alpha479_0_x_locator0);
  gfmult gfm_alpha479_1_x_locator1(10'b1111011111, locator1, alpha479_1_x_locator1);
  gfmult gfm_alpha479_2_x_locator2(10'b1010110011, locator2, alpha479_2_x_locator2);
  gfmult gfm_alpha479_3_x_locator3(10'b1001001110, locator3, alpha479_3_x_locator3);
  gfmult gfm_alpha480_0_x_locator0(10'b0000000001, locator0, alpha480_0_x_locator0);
  gfmult gfm_alpha480_1_x_locator1(10'b1111101011, locator1, alpha480_1_x_locator1);
  gfmult gfm_alpha480_2_x_locator2(10'b1110101010, locator2, alpha480_2_x_locator2);
  gfmult gfm_alpha480_3_x_locator3(10'b1101001111, locator3, alpha480_3_x_locator3);
  gfmult gfm_alpha481_0_x_locator0(10'b0000000001, locator0, alpha481_0_x_locator0);
  gfmult gfm_alpha481_1_x_locator1(10'b1111110001, locator1, alpha481_1_x_locator1);
  gfmult gfm_alpha481_2_x_locator2(10'b1011101110, locator2, alpha481_2_x_locator2);
  gfmult gfm_alpha481_3_x_locator3(10'b1111101110, locator3, alpha481_3_x_locator3);
  gfmult gfm_alpha482_0_x_locator0(10'b0000000001, locator0, alpha482_0_x_locator0);
  gfmult gfm_alpha482_1_x_locator1(10'b1111111100, locator1, alpha482_1_x_locator1);
  gfmult gfm_alpha482_2_x_locator2(10'b1010111111, locator2, alpha482_2_x_locator2);
  gfmult gfm_alpha482_3_x_locator3(10'b1101111011, locator3, alpha482_3_x_locator3);
  gfmult gfm_alpha483_0_x_locator0(10'b0000000001, locator0, alpha483_0_x_locator0);
  gfmult gfm_alpha483_1_x_locator1(10'b0111111110, locator1, alpha483_1_x_locator1);
  gfmult gfm_alpha483_2_x_locator2(10'b1110101001, locator2, alpha483_2_x_locator2);
  gfmult gfm_alpha483_3_x_locator3(10'b0111101100, locator3, alpha483_3_x_locator3);
  gfmult gfm_alpha484_0_x_locator0(10'b0000000001, locator0, alpha484_0_x_locator0);
  gfmult gfm_alpha484_1_x_locator1(10'b0011111111, locator1, alpha484_1_x_locator1);
  gfmult gfm_alpha484_2_x_locator2(10'b0111101000, locator2, alpha484_2_x_locator2);
  gfmult gfm_alpha484_3_x_locator3(10'b1000111001, locator3, alpha484_3_x_locator3);
  gfmult gfm_alpha485_0_x_locator0(10'b0000000001, locator0, alpha485_0_x_locator0);
  gfmult gfm_alpha485_1_x_locator1(10'b1001111011, locator1, alpha485_1_x_locator1);
  gfmult gfm_alpha485_2_x_locator2(10'b0001111010, locator2, alpha485_2_x_locator2);
  gfmult gfm_alpha485_3_x_locator3(10'b0011000110, locator3, alpha485_3_x_locator3);
  gfmult gfm_alpha486_0_x_locator0(10'b0000000001, locator0, alpha486_0_x_locator0);
  gfmult gfm_alpha486_1_x_locator1(10'b1100111001, locator1, alpha486_1_x_locator1);
  gfmult gfm_alpha486_2_x_locator2(10'b1000011010, locator2, alpha486_2_x_locator2);
  gfmult gfm_alpha486_3_x_locator3(10'b1100011110, locator3, alpha486_3_x_locator3);
  gfmult gfm_alpha487_0_x_locator0(10'b0000000001, locator0, alpha487_0_x_locator0);
  gfmult gfm_alpha487_1_x_locator1(10'b1110011000, locator1, alpha487_1_x_locator1);
  gfmult gfm_alpha487_2_x_locator2(10'b1010000010, locator2, alpha487_2_x_locator2);
  gfmult gfm_alpha487_3_x_locator3(10'b1101100101, locator3, alpha487_3_x_locator3);
  gfmult gfm_alpha488_0_x_locator0(10'b0000000001, locator0, alpha488_0_x_locator0);
  gfmult gfm_alpha488_1_x_locator1(10'b0111001100, locator1, alpha488_1_x_locator1);
  gfmult gfm_alpha488_2_x_locator2(10'b1010100100, locator2, alpha488_2_x_locator2);
  gfmult gfm_alpha488_3_x_locator3(10'b1011101001, locator3, alpha488_3_x_locator3);
  gfmult gfm_alpha489_0_x_locator0(10'b0000000001, locator0, alpha489_0_x_locator0);
  gfmult gfm_alpha489_1_x_locator1(10'b0011100110, locator1, alpha489_1_x_locator1);
  gfmult gfm_alpha489_2_x_locator2(10'b0010101001, locator2, alpha489_2_x_locator2);
  gfmult gfm_alpha489_3_x_locator3(10'b0011011100, locator3, alpha489_3_x_locator3);
  gfmult gfm_alpha490_0_x_locator0(10'b0000000001, locator0, alpha490_0_x_locator0);
  gfmult gfm_alpha490_1_x_locator1(10'b0001110011, locator1, alpha490_1_x_locator1);
  gfmult gfm_alpha490_2_x_locator2(10'b0100101000, locator2, alpha490_2_x_locator2);
  gfmult gfm_alpha490_3_x_locator3(10'b1000011111, locator3, alpha490_3_x_locator3);
  gfmult gfm_alpha491_0_x_locator0(10'b0000000001, locator0, alpha491_0_x_locator0);
  gfmult gfm_alpha491_1_x_locator1(10'b1000111101, locator1, alpha491_1_x_locator1);
  gfmult gfm_alpha491_2_x_locator2(10'b0001001010, locator2, alpha491_2_x_locator2);
  gfmult gfm_alpha491_3_x_locator3(10'b1111000100, locator3, alpha491_3_x_locator3);
  gfmult gfm_alpha492_0_x_locator0(10'b0000000001, locator0, alpha492_0_x_locator0);
  gfmult gfm_alpha492_1_x_locator1(10'b1100011010, locator1, alpha492_1_x_locator1);
  gfmult gfm_alpha492_2_x_locator2(10'b1000010110, locator2, alpha492_2_x_locator2);
  gfmult gfm_alpha492_3_x_locator3(10'b1001111100, locator3, alpha492_3_x_locator3);
  gfmult gfm_alpha493_0_x_locator0(10'b0000000001, locator0, alpha493_0_x_locator0);
  gfmult gfm_alpha493_1_x_locator1(10'b0110001101, locator1, alpha493_1_x_locator1);
  gfmult gfm_alpha493_2_x_locator2(10'b1010000001, locator2, alpha493_2_x_locator2);
  gfmult gfm_alpha493_3_x_locator3(10'b1001001011, locator3, alpha493_3_x_locator3);
  gfmult gfm_alpha494_0_x_locator0(10'b0000000001, locator0, alpha494_0_x_locator0);
  gfmult gfm_alpha494_1_x_locator1(10'b1011000010, locator1, alpha494_1_x_locator1);
  gfmult gfm_alpha494_2_x_locator2(10'b0110100010, locator2, alpha494_2_x_locator2);
  gfmult gfm_alpha494_3_x_locator3(10'b0111001010, locator3, alpha494_3_x_locator3);
  gfmult gfm_alpha495_0_x_locator0(10'b0000000001, locator0, alpha495_0_x_locator0);
  gfmult gfm_alpha495_1_x_locator1(10'b0101100001, locator1, alpha495_1_x_locator1);
  gfmult gfm_alpha495_2_x_locator2(10'b1001101100, locator2, alpha495_2_x_locator2);
  gfmult gfm_alpha495_3_x_locator3(10'b0100111011, locator3, alpha495_3_x_locator3);
  gfmult gfm_alpha496_0_x_locator0(10'b0000000001, locator0, alpha496_0_x_locator0);
  gfmult gfm_alpha496_1_x_locator1(10'b1010110100, locator1, alpha496_1_x_locator1);
  gfmult gfm_alpha496_2_x_locator2(10'b0010011011, locator2, alpha496_2_x_locator2);
  gfmult gfm_alpha496_3_x_locator3(10'b0110100100, locator3, alpha496_3_x_locator3);
  gfmult gfm_alpha497_0_x_locator0(10'b0000000001, locator0, alpha497_0_x_locator0);
  gfmult gfm_alpha497_1_x_locator1(10'b0101011010, locator1, alpha497_1_x_locator1);
  gfmult gfm_alpha497_2_x_locator2(10'b1100100000, locator2, alpha497_2_x_locator2);
  gfmult gfm_alpha497_3_x_locator3(10'b1000110000, locator3, alpha497_3_x_locator3);
  gfmult gfm_alpha498_0_x_locator0(10'b0000000001, locator0, alpha498_0_x_locator0);
  gfmult gfm_alpha498_1_x_locator1(10'b0010101101, locator1, alpha498_1_x_locator1);
  gfmult gfm_alpha498_2_x_locator2(10'b0011001000, locator2, alpha498_2_x_locator2);
  gfmult gfm_alpha498_3_x_locator3(10'b0001000110, locator3, alpha498_3_x_locator3);
  gfmult gfm_alpha499_0_x_locator0(10'b0000000001, locator0, alpha499_0_x_locator0);
  gfmult gfm_alpha499_1_x_locator1(10'b1001010010, locator1, alpha499_1_x_locator1);
  gfmult gfm_alpha499_2_x_locator2(10'b0000110010, locator2, alpha499_2_x_locator2);
  gfmult gfm_alpha499_3_x_locator3(10'b1100001110, locator3, alpha499_3_x_locator3);
  gfmult gfm_alpha500_0_x_locator0(10'b0000000001, locator0, alpha500_0_x_locator0);
  gfmult gfm_alpha500_1_x_locator1(10'b0100101001, locator1, alpha500_1_x_locator1);
  gfmult gfm_alpha500_2_x_locator2(10'b1000001000, locator2, alpha500_2_x_locator2);
  gfmult gfm_alpha500_3_x_locator3(10'b1101100111, locator3, alpha500_3_x_locator3);
  gfmult gfm_alpha501_0_x_locator0(10'b0000000001, locator0, alpha501_0_x_locator0);
  gfmult gfm_alpha501_1_x_locator1(10'b1010010000, locator1, alpha501_1_x_locator1);
  gfmult gfm_alpha501_2_x_locator2(10'b0010000010, locator2, alpha501_2_x_locator2);
  gfmult gfm_alpha501_3_x_locator3(10'b1111101011, locator3, alpha501_3_x_locator3);
  gfmult gfm_alpha502_0_x_locator0(10'b0000000001, locator0, alpha502_0_x_locator0);
  gfmult gfm_alpha502_1_x_locator1(10'b0101001000, locator1, alpha502_1_x_locator1);
  gfmult gfm_alpha502_2_x_locator2(10'b1000100100, locator2, alpha502_2_x_locator2);
  gfmult gfm_alpha502_3_x_locator3(10'b0111111110, locator3, alpha502_3_x_locator3);
  gfmult gfm_alpha503_0_x_locator0(10'b0000000001, locator0, alpha503_0_x_locator0);
  gfmult gfm_alpha503_1_x_locator1(10'b0010100100, locator1, alpha503_1_x_locator1);
  gfmult gfm_alpha503_2_x_locator2(10'b0010001001, locator2, alpha503_2_x_locator2);
  gfmult gfm_alpha503_3_x_locator3(10'b1100111001, locator3, alpha503_3_x_locator3);
  gfmult gfm_alpha504_0_x_locator0(10'b0000000001, locator0, alpha504_0_x_locator0);
  gfmult gfm_alpha504_1_x_locator1(10'b0001010010, locator1, alpha504_1_x_locator1);
  gfmult gfm_alpha504_2_x_locator2(10'b0100100000, locator2, alpha504_2_x_locator2);
  gfmult gfm_alpha504_3_x_locator3(10'b0011100110, locator3, alpha504_3_x_locator3);
  gfmult gfm_alpha505_0_x_locator0(10'b0000000001, locator0, alpha505_0_x_locator0);
  gfmult gfm_alpha505_1_x_locator1(10'b0000101001, locator1, alpha505_1_x_locator1);
  gfmult gfm_alpha505_2_x_locator2(10'b0001001000, locator2, alpha505_2_x_locator2);
  gfmult gfm_alpha505_3_x_locator3(10'b1100011010, locator3, alpha505_3_x_locator3);
  gfmult gfm_alpha506_0_x_locator0(10'b0000000001, locator0, alpha506_0_x_locator0);
  gfmult gfm_alpha506_1_x_locator1(10'b1000010000, locator1, alpha506_1_x_locator1);
  gfmult gfm_alpha506_2_x_locator2(10'b0000010010, locator2, alpha506_2_x_locator2);
  gfmult gfm_alpha506_3_x_locator3(10'b0101100001, locator3, alpha506_3_x_locator3);
  gfmult gfm_alpha507_0_x_locator0(10'b0000000001, locator0, alpha507_0_x_locator0);
  gfmult gfm_alpha507_1_x_locator1(10'b0100001000, locator1, alpha507_1_x_locator1);
  gfmult gfm_alpha507_2_x_locator2(10'b1000000000, locator2, alpha507_2_x_locator2);
  gfmult gfm_alpha507_3_x_locator3(10'b0010101101, locator3, alpha507_3_x_locator3);
  gfmult gfm_alpha508_0_x_locator0(10'b0000000001, locator0, alpha508_0_x_locator0);
  gfmult gfm_alpha508_1_x_locator1(10'b0010000100, locator1, alpha508_1_x_locator1);
  gfmult gfm_alpha508_2_x_locator2(10'b0010000000, locator2, alpha508_2_x_locator2);
  gfmult gfm_alpha508_3_x_locator3(10'b1010010000, locator3, alpha508_3_x_locator3);
  gfmult gfm_alpha509_0_x_locator0(10'b0000000001, locator0, alpha509_0_x_locator0);
  gfmult gfm_alpha509_1_x_locator1(10'b0001000010, locator1, alpha509_1_x_locator1);
  gfmult gfm_alpha509_2_x_locator2(10'b0000100000, locator2, alpha509_2_x_locator2);
  gfmult gfm_alpha509_3_x_locator3(10'b0001010010, locator3, alpha509_3_x_locator3);
  gfmult gfm_alpha510_0_x_locator0(10'b0000000001, locator0, alpha510_0_x_locator0);
  gfmult gfm_alpha510_1_x_locator1(10'b0000100001, locator1, alpha510_1_x_locator1);
  gfmult gfm_alpha510_2_x_locator2(10'b0000001000, locator2, alpha510_2_x_locator2);
  gfmult gfm_alpha510_3_x_locator3(10'b0100001000, locator3, alpha510_3_x_locator3);
  gfmult gfm_alpha511_0_x_locator0(10'b0000000001, locator0, alpha511_0_x_locator0);
  gfmult gfm_alpha511_1_x_locator1(10'b1000010100, locator1, alpha511_1_x_locator1);
  gfmult gfm_alpha511_2_x_locator2(10'b0000000010, locator2, alpha511_2_x_locator2);
  gfmult gfm_alpha511_3_x_locator3(10'b0000100001, locator3, alpha511_3_x_locator3);
  gfmult gfm_alpha512_0_x_locator0(10'b0000000001, locator0, alpha512_0_x_locator0);
  gfmult gfm_alpha512_1_x_locator1(10'b0100001010, locator1, alpha512_1_x_locator1);
  gfmult gfm_alpha512_2_x_locator2(10'b1000000100, locator2, alpha512_2_x_locator2);
  gfmult gfm_alpha512_3_x_locator3(10'b0010000101, locator3, alpha512_3_x_locator3);
  gfmult gfm_alpha513_0_x_locator0(10'b0000000001, locator0, alpha513_0_x_locator0);
  gfmult gfm_alpha513_1_x_locator1(10'b0010000101, locator1, alpha513_1_x_locator1);
  gfmult gfm_alpha513_2_x_locator2(10'b0010000001, locator2, alpha513_2_x_locator2);
  gfmult gfm_alpha513_3_x_locator3(10'b1010010101, locator3, alpha513_3_x_locator3);
  gfmult gfm_alpha514_0_x_locator0(10'b0000000001, locator0, alpha514_0_x_locator0);
  gfmult gfm_alpha514_1_x_locator1(10'b1001000110, locator1, alpha514_1_x_locator1);
  gfmult gfm_alpha514_2_x_locator2(10'b0100100010, locator2, alpha514_2_x_locator2);
  gfmult gfm_alpha514_3_x_locator3(10'b1011010111, locator3, alpha514_3_x_locator3);
  gfmult gfm_alpha515_0_x_locator0(10'b0000000001, locator0, alpha515_0_x_locator0);
  gfmult gfm_alpha515_1_x_locator1(10'b0100100011, locator1, alpha515_1_x_locator1);
  gfmult gfm_alpha515_2_x_locator2(10'b1001001100, locator2, alpha515_2_x_locator2);
  gfmult gfm_alpha515_3_x_locator3(10'b1111011101, locator3, alpha515_3_x_locator3);
  gfmult gfm_alpha516_0_x_locator0(10'b0000000001, locator0, alpha516_0_x_locator0);
  gfmult gfm_alpha516_1_x_locator1(10'b1010010101, locator1, alpha516_1_x_locator1);
  gfmult gfm_alpha516_2_x_locator2(10'b0010010011, locator2, alpha516_2_x_locator2);
  gfmult gfm_alpha516_3_x_locator3(10'b1011111110, locator3, alpha516_3_x_locator3);
  gfmult gfm_alpha517_0_x_locator0(10'b0000000001, locator0, alpha517_0_x_locator0);
  gfmult gfm_alpha517_1_x_locator1(10'b1101001110, locator1, alpha517_1_x_locator1);
  gfmult gfm_alpha517_2_x_locator2(10'b1100100010, locator2, alpha517_2_x_locator2);
  gfmult gfm_alpha517_3_x_locator3(10'b1101011001, locator3, alpha517_3_x_locator3);
  gfmult gfm_alpha518_0_x_locator0(10'b0000000001, locator0, alpha518_0_x_locator0);
  gfmult gfm_alpha518_1_x_locator1(10'b0110100111, locator1, alpha518_1_x_locator1);
  gfmult gfm_alpha518_2_x_locator2(10'b1011001100, locator2, alpha518_2_x_locator2);
  gfmult gfm_alpha518_3_x_locator3(10'b0011101010, locator3, alpha518_3_x_locator3);
  gfmult gfm_alpha519_0_x_locator0(10'b0000000001, locator0, alpha519_0_x_locator0);
  gfmult gfm_alpha519_1_x_locator1(10'b1011010111, locator1, alpha519_1_x_locator1);
  gfmult gfm_alpha519_2_x_locator2(10'b0010110011, locator2, alpha519_2_x_locator2);
  gfmult gfm_alpha519_3_x_locator3(10'b0100011111, locator3, alpha519_3_x_locator3);
  gfmult gfm_alpha520_0_x_locator0(10'b0000000001, locator0, alpha520_0_x_locator0);
  gfmult gfm_alpha520_1_x_locator1(10'b1101101111, locator1, alpha520_1_x_locator1);
  gfmult gfm_alpha520_2_x_locator2(10'b1100101010, locator2, alpha520_2_x_locator2);
  gfmult gfm_alpha520_3_x_locator3(10'b1110100100, locator3, alpha520_3_x_locator3);
  gfmult gfm_alpha521_0_x_locator0(10'b0000000001, locator0, alpha521_0_x_locator0);
  gfmult gfm_alpha521_1_x_locator1(10'b1110110011, locator1, alpha521_1_x_locator1);
  gfmult gfm_alpha521_2_x_locator2(10'b1011001110, locator2, alpha521_2_x_locator2);
  gfmult gfm_alpha521_3_x_locator3(10'b1001110000, locator3, alpha521_3_x_locator3);
  gfmult gfm_alpha522_0_x_locator0(10'b0000000001, locator0, alpha522_0_x_locator0);
  gfmult gfm_alpha522_1_x_locator1(10'b1111011101, locator1, alpha522_1_x_locator1);
  gfmult gfm_alpha522_2_x_locator2(10'b1010110111, locator2, alpha522_2_x_locator2);
  gfmult gfm_alpha522_3_x_locator3(10'b0001001110, locator3, alpha522_3_x_locator3);
  gfmult gfm_alpha523_0_x_locator0(10'b0000000001, locator0, alpha523_0_x_locator0);
  gfmult gfm_alpha523_1_x_locator1(10'b1111101010, locator1, alpha523_1_x_locator1);
  gfmult gfm_alpha523_2_x_locator2(10'b1110101011, locator2, alpha523_2_x_locator2);
  gfmult gfm_alpha523_3_x_locator3(10'b1100001111, locator3, alpha523_3_x_locator3);
  gfmult gfm_alpha524_0_x_locator0(10'b0000000001, locator0, alpha524_0_x_locator0);
  gfmult gfm_alpha524_1_x_locator1(10'b0111110101, locator1, alpha524_1_x_locator1);
  gfmult gfm_alpha524_2_x_locator2(10'b1111101100, locator2, alpha524_2_x_locator2);
  gfmult gfm_alpha524_3_x_locator3(10'b1111100110, locator3, alpha524_3_x_locator3);
  gfmult gfm_alpha525_0_x_locator0(10'b0000000001, locator0, alpha525_0_x_locator0);
  gfmult gfm_alpha525_1_x_locator1(10'b1011111110, locator1, alpha525_1_x_locator1);
  gfmult gfm_alpha525_2_x_locator2(10'b0011111011, locator2, alpha525_2_x_locator2);
  gfmult gfm_alpha525_3_x_locator3(10'b1101111010, locator3, alpha525_3_x_locator3);
  gfmult gfm_alpha526_0_x_locator0(10'b0000000001, locator0, alpha526_0_x_locator0);
  gfmult gfm_alpha526_1_x_locator1(10'b0101111111, locator1, alpha526_1_x_locator1);
  gfmult gfm_alpha526_2_x_locator2(10'b1100111000, locator2, alpha526_2_x_locator2);
  gfmult gfm_alpha526_3_x_locator3(10'b0101101101, locator3, alpha526_3_x_locator3);
  gfmult gfm_alpha527_0_x_locator0(10'b0000000001, locator0, alpha527_0_x_locator0);
  gfmult gfm_alpha527_1_x_locator1(10'b1010111011, locator1, alpha527_1_x_locator1);
  gfmult gfm_alpha527_2_x_locator2(10'b0011001110, locator2, alpha527_2_x_locator2);
  gfmult gfm_alpha527_3_x_locator3(10'b1010101000, locator3, alpha527_3_x_locator3);
  gfmult gfm_alpha528_0_x_locator0(10'b0000000001, locator0, alpha528_0_x_locator0);
  gfmult gfm_alpha528_1_x_locator1(10'b1101011001, locator1, alpha528_1_x_locator1);
  gfmult gfm_alpha528_2_x_locator2(10'b1000110111, locator2, alpha528_2_x_locator2);
  gfmult gfm_alpha528_3_x_locator3(10'b0001010101, locator3, alpha528_3_x_locator3);
  gfmult gfm_alpha529_0_x_locator0(10'b0000000001, locator0, alpha529_0_x_locator0);
  gfmult gfm_alpha529_1_x_locator1(10'b1110101000, locator1, alpha529_1_x_locator1);
  gfmult gfm_alpha529_2_x_locator2(10'b1110001011, locator2, alpha529_2_x_locator2);
  gfmult gfm_alpha529_3_x_locator3(10'b1010001111, locator3, alpha529_3_x_locator3);
  gfmult gfm_alpha530_0_x_locator0(10'b0000000001, locator0, alpha530_0_x_locator0);
  gfmult gfm_alpha530_1_x_locator1(10'b0111010100, locator1, alpha530_1_x_locator1);
  gfmult gfm_alpha530_2_x_locator2(10'b1111100100, locator2, alpha530_2_x_locator2);
  gfmult gfm_alpha530_3_x_locator3(10'b1111010110, locator3, alpha530_3_x_locator3);
  gfmult gfm_alpha531_0_x_locator0(10'b0000000001, locator0, alpha531_0_x_locator0);
  gfmult gfm_alpha531_1_x_locator1(10'b0011101010, locator1, alpha531_1_x_locator1);
  gfmult gfm_alpha531_2_x_locator2(10'b0011111001, locator2, alpha531_2_x_locator2);
  gfmult gfm_alpha531_3_x_locator3(10'b1101111100, locator3, alpha531_3_x_locator3);
  gfmult gfm_alpha532_0_x_locator0(10'b0000000001, locator0, alpha532_0_x_locator0);
  gfmult gfm_alpha532_1_x_locator1(10'b0001110101, locator1, alpha532_1_x_locator1);
  gfmult gfm_alpha532_2_x_locator2(10'b0100111100, locator2, alpha532_2_x_locator2);
  gfmult gfm_alpha532_3_x_locator3(10'b1001101011, locator3, alpha532_3_x_locator3);
  gfmult gfm_alpha533_0_x_locator0(10'b0000000001, locator0, alpha533_0_x_locator0);
  gfmult gfm_alpha533_1_x_locator1(10'b1000111110, locator1, alpha533_1_x_locator1);
  gfmult gfm_alpha533_2_x_locator2(10'b0001001111, locator2, alpha533_2_x_locator2);
  gfmult gfm_alpha533_3_x_locator3(10'b0111001110, locator3, alpha533_3_x_locator3);
  gfmult gfm_alpha534_0_x_locator0(10'b0000000001, locator0, alpha534_0_x_locator0);
  gfmult gfm_alpha534_1_x_locator1(10'b0100011111, locator1, alpha534_1_x_locator1);
  gfmult gfm_alpha534_2_x_locator2(10'b1100010101, locator2, alpha534_2_x_locator2);
  gfmult gfm_alpha534_3_x_locator3(10'b1100111111, locator3, alpha534_3_x_locator3);
  gfmult gfm_alpha535_0_x_locator0(10'b0000000001, locator0, alpha535_0_x_locator0);
  gfmult gfm_alpha535_1_x_locator1(10'b1010001011, locator1, alpha535_1_x_locator1);
  gfmult gfm_alpha535_2_x_locator2(10'b0111000111, locator2, alpha535_2_x_locator2);
  gfmult gfm_alpha535_3_x_locator3(10'b1111100000, locator3, alpha535_3_x_locator3);
  gfmult gfm_alpha536_0_x_locator0(10'b0000000001, locator0, alpha536_0_x_locator0);
  gfmult gfm_alpha536_1_x_locator1(10'b1101000001, locator1, alpha536_1_x_locator1);
  gfmult gfm_alpha536_2_x_locator2(10'b1101110111, locator2, alpha536_2_x_locator2);
  gfmult gfm_alpha536_3_x_locator3(10'b0001111100, locator3, alpha536_3_x_locator3);
  gfmult gfm_alpha537_0_x_locator0(10'b0000000001, locator0, alpha537_0_x_locator0);
  gfmult gfm_alpha537_1_x_locator1(10'b1110100100, locator1, alpha537_1_x_locator1);
  gfmult gfm_alpha537_2_x_locator2(10'b1111011011, locator2, alpha537_2_x_locator2);
  gfmult gfm_alpha537_3_x_locator3(10'b1000001011, locator3, alpha537_3_x_locator3);
  gfmult gfm_alpha538_0_x_locator0(10'b0000000001, locator0, alpha538_0_x_locator0);
  gfmult gfm_alpha538_1_x_locator1(10'b0111010010, locator1, alpha538_1_x_locator1);
  gfmult gfm_alpha538_2_x_locator2(10'b1111110000, locator2, alpha538_2_x_locator2);
  gfmult gfm_alpha538_3_x_locator3(10'b0111000010, locator3, alpha538_3_x_locator3);
  gfmult gfm_alpha539_0_x_locator0(10'b0000000001, locator0, alpha539_0_x_locator0);
  gfmult gfm_alpha539_1_x_locator1(10'b0011101001, locator1, alpha539_1_x_locator1);
  gfmult gfm_alpha539_2_x_locator2(10'b0011111100, locator2, alpha539_2_x_locator2);
  gfmult gfm_alpha539_3_x_locator3(10'b0100111010, locator3, alpha539_3_x_locator3);
  gfmult gfm_alpha540_0_x_locator0(10'b0000000001, locator0, alpha540_0_x_locator0);
  gfmult gfm_alpha540_1_x_locator1(10'b1001110000, locator1, alpha540_1_x_locator1);
  gfmult gfm_alpha540_2_x_locator2(10'b0000111111, locator2, alpha540_2_x_locator2);
  gfmult gfm_alpha540_3_x_locator3(10'b0100100101, locator3, alpha540_3_x_locator3);
  gfmult gfm_alpha541_0_x_locator0(10'b0000000001, locator0, alpha541_0_x_locator0);
  gfmult gfm_alpha541_1_x_locator1(10'b0100111000, locator1, alpha541_1_x_locator1);
  gfmult gfm_alpha541_2_x_locator2(10'b1100001001, locator2, alpha541_2_x_locator2);
  gfmult gfm_alpha541_3_x_locator3(10'b1010100001, locator3, alpha541_3_x_locator3);

  assign codeword = received ^ error;
  assign error = {(~| (alpha541_0_x_locator0 ^ alpha541_1_x_locator1 ^ alpha541_2_x_locator2 ^ alpha541_3_x_locator3)), 
  (~| (alpha540_0_x_locator0 ^ alpha540_1_x_locator1 ^ alpha540_2_x_locator2 ^ alpha540_3_x_locator3)), 
  (~| (alpha539_0_x_locator0 ^ alpha539_1_x_locator1 ^ alpha539_2_x_locator2 ^ alpha539_3_x_locator3)), 
  (~| (alpha538_0_x_locator0 ^ alpha538_1_x_locator1 ^ alpha538_2_x_locator2 ^ alpha538_3_x_locator3)), 
  (~| (alpha537_0_x_locator0 ^ alpha537_1_x_locator1 ^ alpha537_2_x_locator2 ^ alpha537_3_x_locator3)), 
  (~| (alpha536_0_x_locator0 ^ alpha536_1_x_locator1 ^ alpha536_2_x_locator2 ^ alpha536_3_x_locator3)), 
  (~| (alpha535_0_x_locator0 ^ alpha535_1_x_locator1 ^ alpha535_2_x_locator2 ^ alpha535_3_x_locator3)), 
  (~| (alpha534_0_x_locator0 ^ alpha534_1_x_locator1 ^ alpha534_2_x_locator2 ^ alpha534_3_x_locator3)), 
  (~| (alpha533_0_x_locator0 ^ alpha533_1_x_locator1 ^ alpha533_2_x_locator2 ^ alpha533_3_x_locator3)), (~| (alpha532_0_x_locator0 ^ alpha532_1_x_locator1 ^ alpha532_2_x_locator2 ^ alpha532_3_x_locator3)), (~| (alpha531_0_x_locator0 ^ alpha531_1_x_locator1 ^ alpha531_2_x_locator2 ^ alpha531_3_x_locator3)), (~| (alpha530_0_x_locator0 ^ alpha530_1_x_locator1 ^ alpha530_2_x_locator2 ^ alpha530_3_x_locator3)), (~| (alpha529_0_x_locator0 ^ alpha529_1_x_locator1 ^ alpha529_2_x_locator2 ^ alpha529_3_x_locator3)), (~| (alpha528_0_x_locator0 ^ alpha528_1_x_locator1 ^ alpha528_2_x_locator2 ^ alpha528_3_x_locator3)), (~| (alpha527_0_x_locator0 ^ alpha527_1_x_locator1 ^ alpha527_2_x_locator2 ^ alpha527_3_x_locator3)), (~| (alpha526_0_x_locator0 ^ alpha526_1_x_locator1 ^ alpha526_2_x_locator2 ^ alpha526_3_x_locator3)), (~| (alpha525_0_x_locator0 ^ alpha525_1_x_locator1 ^ alpha525_2_x_locator2 ^ alpha525_3_x_locator3)), (~| (alpha524_0_x_locator0 ^ alpha524_1_x_locator1 ^ alpha524_2_x_locator2 ^ alpha524_3_x_locator3)), (~| (alpha523_0_x_locator0 ^ alpha523_1_x_locator1 ^ alpha523_2_x_locator2 ^ alpha523_3_x_locator3)), (~| (alpha522_0_x_locator0 ^ alpha522_1_x_locator1 ^ alpha522_2_x_locator2 ^ alpha522_3_x_locator3)), (~| (alpha521_0_x_locator0 ^ alpha521_1_x_locator1 ^ alpha521_2_x_locator2 ^ alpha521_3_x_locator3)), (~| (alpha520_0_x_locator0 ^ alpha520_1_x_locator1 ^ alpha520_2_x_locator2 ^ alpha520_3_x_locator3)), (~| (alpha519_0_x_locator0 ^ alpha519_1_x_locator1 ^ alpha519_2_x_locator2 ^ alpha519_3_x_locator3)), (~| (alpha518_0_x_locator0 ^ alpha518_1_x_locator1 ^ alpha518_2_x_locator2 ^ alpha518_3_x_locator3)), (~| (alpha517_0_x_locator0 ^ alpha517_1_x_locator1 ^ alpha517_2_x_locator2 ^ alpha517_3_x_locator3)), (~| (alpha516_0_x_locator0 ^ alpha516_1_x_locator1 ^ alpha516_2_x_locator2 ^ alpha516_3_x_locator3)), (~| (alpha515_0_x_locator0 ^ alpha515_1_x_locator1 ^ alpha515_2_x_locator2 ^ alpha515_3_x_locator3)), (~| (alpha514_0_x_locator0 ^ alpha514_1_x_locator1 ^ alpha514_2_x_locator2 ^ alpha514_3_x_locator3)), (~| (alpha513_0_x_locator0 ^ alpha513_1_x_locator1 ^ alpha513_2_x_locator2 ^ alpha513_3_x_locator3)), (~| (alpha512_0_x_locator0 ^ alpha512_1_x_locator1 ^ alpha512_2_x_locator2 ^ alpha512_3_x_locator3)), (~| (alpha511_0_x_locator0 ^ alpha511_1_x_locator1 ^ alpha511_2_x_locator2 ^ alpha511_3_x_locator3)), (~| (alpha510_0_x_locator0 ^ alpha510_1_x_locator1 ^ alpha510_2_x_locator2 ^ alpha510_3_x_locator3)), (~| (alpha509_0_x_locator0 ^ alpha509_1_x_locator1 ^ alpha509_2_x_locator2 ^ alpha509_3_x_locator3)), (~| (alpha508_0_x_locator0 ^ alpha508_1_x_locator1 ^ alpha508_2_x_locator2 ^ alpha508_3_x_locator3)), (~| (alpha507_0_x_locator0 ^ alpha507_1_x_locator1 ^ alpha507_2_x_locator2 ^ alpha507_3_x_locator3)), (~| (alpha506_0_x_locator0 ^ alpha506_1_x_locator1 ^ alpha506_2_x_locator2 ^ alpha506_3_x_locator3)), (~| (alpha505_0_x_locator0 ^ alpha505_1_x_locator1 ^ alpha505_2_x_locator2 ^ alpha505_3_x_locator3)), (~| (alpha504_0_x_locator0 ^ alpha504_1_x_locator1 ^ alpha504_2_x_locator2 ^ alpha504_3_x_locator3)), (~| (alpha503_0_x_locator0 ^ alpha503_1_x_locator1 ^ alpha503_2_x_locator2 ^ alpha503_3_x_locator3)), (~| (alpha502_0_x_locator0 ^ alpha502_1_x_locator1 ^ alpha502_2_x_locator2 ^ alpha502_3_x_locator3)), (~| (alpha501_0_x_locator0 ^ alpha501_1_x_locator1 ^ alpha501_2_x_locator2 ^ alpha501_3_x_locator3)), (~| (alpha500_0_x_locator0 ^ alpha500_1_x_locator1 ^ alpha500_2_x_locator2 ^ alpha500_3_x_locator3)), (~| (alpha499_0_x_locator0 ^ alpha499_1_x_locator1 ^ alpha499_2_x_locator2 ^ alpha499_3_x_locator3)), (~| (alpha498_0_x_locator0 ^ alpha498_1_x_locator1 ^ alpha498_2_x_locator2 ^ alpha498_3_x_locator3)), (~| (alpha497_0_x_locator0 ^ alpha497_1_x_locator1 ^ alpha497_2_x_locator2 ^ alpha497_3_x_locator3)), (~| (alpha496_0_x_locator0 ^ alpha496_1_x_locator1 ^ alpha496_2_x_locator2 ^ alpha496_3_x_locator3)), (~| (alpha495_0_x_locator0 ^ alpha495_1_x_locator1 ^ alpha495_2_x_locator2 ^ alpha495_3_x_locator3)), (~| (alpha494_0_x_locator0 ^ alpha494_1_x_locator1 ^ alpha494_2_x_locator2 ^ alpha494_3_x_locator3)), (~| (alpha493_0_x_locator0 ^ alpha493_1_x_locator1 ^ alpha493_2_x_locator2 ^ alpha493_3_x_locator3)), (~| (alpha492_0_x_locator0 ^ alpha492_1_x_locator1 ^ alpha492_2_x_locator2 ^ alpha492_3_x_locator3)), (~| (alpha491_0_x_locator0 ^ alpha491_1_x_locator1 ^ alpha491_2_x_locator2 ^ alpha491_3_x_locator3)), (~| (alpha490_0_x_locator0 ^ alpha490_1_x_locator1 ^ alpha490_2_x_locator2 ^ alpha490_3_x_locator3)), (~| (alpha489_0_x_locator0 ^ alpha489_1_x_locator1 ^ alpha489_2_x_locator2 ^ alpha489_3_x_locator3)), (~| (alpha488_0_x_locator0 ^ alpha488_1_x_locator1 ^ alpha488_2_x_locator2 ^ alpha488_3_x_locator3)), (~| (alpha487_0_x_locator0 ^ alpha487_1_x_locator1 ^ alpha487_2_x_locator2 ^ alpha487_3_x_locator3)), (~| (alpha486_0_x_locator0 ^ alpha486_1_x_locator1 ^ alpha486_2_x_locator2 ^ alpha486_3_x_locator3)), (~| (alpha485_0_x_locator0 ^ alpha485_1_x_locator1 ^ alpha485_2_x_locator2 ^ alpha485_3_x_locator3)), (~| (alpha484_0_x_locator0 ^ alpha484_1_x_locator1 ^ alpha484_2_x_locator2 ^ alpha484_3_x_locator3)), (~| (alpha483_0_x_locator0 ^ alpha483_1_x_locator1 ^ alpha483_2_x_locator2 ^ alpha483_3_x_locator3)), (~| (alpha482_0_x_locator0 ^ alpha482_1_x_locator1 ^ alpha482_2_x_locator2 ^ alpha482_3_x_locator3)), (~| (alpha481_0_x_locator0 ^ alpha481_1_x_locator1 ^ alpha481_2_x_locator2 ^ alpha481_3_x_locator3)), (~| (alpha480_0_x_locator0 ^ alpha480_1_x_locator1 ^ alpha480_2_x_locator2 ^ alpha480_3_x_locator3)), (~| (alpha479_0_x_locator0 ^ alpha479_1_x_locator1 ^ alpha479_2_x_locator2 ^ alpha479_3_x_locator3)), (~| (alpha478_0_x_locator0 ^ alpha478_1_x_locator1 ^ alpha478_2_x_locator2 ^ alpha478_3_x_locator3)), (~| (alpha477_0_x_locator0 ^ alpha477_1_x_locator1 ^ alpha477_2_x_locator2 ^ alpha477_3_x_locator3)), (~| (alpha476_0_x_locator0 ^ alpha476_1_x_locator1 ^ alpha476_2_x_locator2 ^ alpha476_3_x_locator3)), (~| (alpha475_0_x_locator0 ^ alpha475_1_x_locator1 ^ alpha475_2_x_locator2 ^ alpha475_3_x_locator3)), (~| (alpha474_0_x_locator0 ^ alpha474_1_x_locator1 ^ alpha474_2_x_locator2 ^ alpha474_3_x_locator3)), (~| (alpha473_0_x_locator0 ^ alpha473_1_x_locator1 ^ alpha473_2_x_locator2 ^ alpha473_3_x_locator3)), (~| (alpha472_0_x_locator0 ^ alpha472_1_x_locator1 ^ alpha472_2_x_locator2 ^ alpha472_3_x_locator3)), (~| (alpha471_0_x_locator0 ^ alpha471_1_x_locator1 ^ alpha471_2_x_locator2 ^ alpha471_3_x_locator3)), (~| (alpha470_0_x_locator0 ^ alpha470_1_x_locator1 ^ alpha470_2_x_locator2 ^ alpha470_3_x_locator3)), (~| (alpha469_0_x_locator0 ^ alpha469_1_x_locator1 ^ alpha469_2_x_locator2 ^ alpha469_3_x_locator3)), (~| (alpha468_0_x_locator0 ^ alpha468_1_x_locator1 ^ alpha468_2_x_locator2 ^ alpha468_3_x_locator3)), (~| (alpha467_0_x_locator0 ^ alpha467_1_x_locator1 ^ alpha467_2_x_locator2 ^ alpha467_3_x_locator3)), (~| (alpha466_0_x_locator0 ^ alpha466_1_x_locator1 ^ alpha466_2_x_locator2 ^ alpha466_3_x_locator3)), (~| (alpha465_0_x_locator0 ^ alpha465_1_x_locator1 ^ alpha465_2_x_locator2 ^ alpha465_3_x_locator3)), (~| (alpha464_0_x_locator0 ^ alpha464_1_x_locator1 ^ alpha464_2_x_locator2 ^ alpha464_3_x_locator3)), (~| (alpha463_0_x_locator0 ^ alpha463_1_x_locator1 ^ alpha463_2_x_locator2 ^ alpha463_3_x_locator3)), (~| (alpha462_0_x_locator0 ^ alpha462_1_x_locator1 ^ alpha462_2_x_locator2 ^ alpha462_3_x_locator3)), (~| (alpha461_0_x_locator0 ^ alpha461_1_x_locator1 ^ alpha461_2_x_locator2 ^ alpha461_3_x_locator3)), (~| (alpha460_0_x_locator0 ^ alpha460_1_x_locator1 ^ alpha460_2_x_locator2 ^ alpha460_3_x_locator3)), (~| (alpha459_0_x_locator0 ^ alpha459_1_x_locator1 ^ alpha459_2_x_locator2 ^ alpha459_3_x_locator3)), (~| (alpha458_0_x_locator0 ^ alpha458_1_x_locator1 ^ alpha458_2_x_locator2 ^ alpha458_3_x_locator3)), (~| (alpha457_0_x_locator0 ^ alpha457_1_x_locator1 ^ alpha457_2_x_locator2 ^ alpha457_3_x_locator3)), (~| (alpha456_0_x_locator0 ^ alpha456_1_x_locator1 ^ alpha456_2_x_locator2 ^ alpha456_3_x_locator3)), (~| (alpha455_0_x_locator0 ^ alpha455_1_x_locator1 ^ alpha455_2_x_locator2 ^ alpha455_3_x_locator3)), (~| (alpha454_0_x_locator0 ^ alpha454_1_x_locator1 ^ alpha454_2_x_locator2 ^ alpha454_3_x_locator3)), (~| (alpha453_0_x_locator0 ^ alpha453_1_x_locator1 ^ alpha453_2_x_locator2 ^ alpha453_3_x_locator3)), (~| (alpha452_0_x_locator0 ^ alpha452_1_x_locator1 ^ alpha452_2_x_locator2 ^ alpha452_3_x_locator3)), (~| (alpha451_0_x_locator0 ^ alpha451_1_x_locator1 ^ alpha451_2_x_locator2 ^ alpha451_3_x_locator3)), (~| (alpha450_0_x_locator0 ^ alpha450_1_x_locator1 ^ alpha450_2_x_locator2 ^ alpha450_3_x_locator3)), (~| (alpha449_0_x_locator0 ^ alpha449_1_x_locator1 ^ alpha449_2_x_locator2 ^ alpha449_3_x_locator3)), (~| (alpha448_0_x_locator0 ^ alpha448_1_x_locator1 ^ alpha448_2_x_locator2 ^ alpha448_3_x_locator3)), (~| (alpha447_0_x_locator0 ^ alpha447_1_x_locator1 ^ alpha447_2_x_locator2 ^ alpha447_3_x_locator3)), (~| (alpha446_0_x_locator0 ^ alpha446_1_x_locator1 ^ alpha446_2_x_locator2 ^ alpha446_3_x_locator3)), (~| (alpha445_0_x_locator0 ^ alpha445_1_x_locator1 ^ alpha445_2_x_locator2 ^ alpha445_3_x_locator3)), (~| (alpha444_0_x_locator0 ^ alpha444_1_x_locator1 ^ alpha444_2_x_locator2 ^ alpha444_3_x_locator3)), (~| (alpha443_0_x_locator0 ^ alpha443_1_x_locator1 ^ alpha443_2_x_locator2 ^ alpha443_3_x_locator3)), (~| (alpha442_0_x_locator0 ^ alpha442_1_x_locator1 ^ alpha442_2_x_locator2 ^ alpha442_3_x_locator3)), (~| (alpha441_0_x_locator0 ^ alpha441_1_x_locator1 ^ alpha441_2_x_locator2 ^ alpha441_3_x_locator3)), (~| (alpha440_0_x_locator0 ^ alpha440_1_x_locator1 ^ alpha440_2_x_locator2 ^ alpha440_3_x_locator3)), (~| (alpha439_0_x_locator0 ^ alpha439_1_x_locator1 ^ alpha439_2_x_locator2 ^ alpha439_3_x_locator3)), (~| (alpha438_0_x_locator0 ^ alpha438_1_x_locator1 ^ alpha438_2_x_locator2 ^ alpha438_3_x_locator3)), (~| (alpha437_0_x_locator0 ^ alpha437_1_x_locator1 ^ alpha437_2_x_locator2 ^ alpha437_3_x_locator3)), (~| (alpha436_0_x_locator0 ^ alpha436_1_x_locator1 ^ alpha436_2_x_locator2 ^ alpha436_3_x_locator3)), (~| (alpha435_0_x_locator0 ^ alpha435_1_x_locator1 ^ alpha435_2_x_locator2 ^ alpha435_3_x_locator3)), (~| (alpha434_0_x_locator0 ^ alpha434_1_x_locator1 ^ alpha434_2_x_locator2 ^ alpha434_3_x_locator3)), (~| (alpha433_0_x_locator0 ^ alpha433_1_x_locator1 ^ alpha433_2_x_locator2 ^ alpha433_3_x_locator3)), (~| (alpha432_0_x_locator0 ^ alpha432_1_x_locator1 ^ alpha432_2_x_locator2 ^ alpha432_3_x_locator3)), (~| (alpha431_0_x_locator0 ^ alpha431_1_x_locator1 ^ alpha431_2_x_locator2 ^ alpha431_3_x_locator3)), (~| (alpha430_0_x_locator0 ^ alpha430_1_x_locator1 ^ alpha430_2_x_locator2 ^ alpha430_3_x_locator3)), (~| (alpha429_0_x_locator0 ^ alpha429_1_x_locator1 ^ alpha429_2_x_locator2 ^ alpha429_3_x_locator3)), (~| (alpha428_0_x_locator0 ^ alpha428_1_x_locator1 ^ alpha428_2_x_locator2 ^ alpha428_3_x_locator3)), (~| (alpha427_0_x_locator0 ^ alpha427_1_x_locator1 ^ alpha427_2_x_locator2 ^ alpha427_3_x_locator3)), (~| (alpha426_0_x_locator0 ^ alpha426_1_x_locator1 ^ alpha426_2_x_locator2 ^ alpha426_3_x_locator3)), (~| (alpha425_0_x_locator0 ^ alpha425_1_x_locator1 ^ alpha425_2_x_locator2 ^ alpha425_3_x_locator3)), (~| (alpha424_0_x_locator0 ^ alpha424_1_x_locator1 ^ alpha424_2_x_locator2 ^ alpha424_3_x_locator3)), (~| (alpha423_0_x_locator0 ^ alpha423_1_x_locator1 ^ alpha423_2_x_locator2 ^ alpha423_3_x_locator3)), (~| (alpha422_0_x_locator0 ^ alpha422_1_x_locator1 ^ alpha422_2_x_locator2 ^ alpha422_3_x_locator3)), (~| (alpha421_0_x_locator0 ^ alpha421_1_x_locator1 ^ alpha421_2_x_locator2 ^ alpha421_3_x_locator3)), (~| (alpha420_0_x_locator0 ^ alpha420_1_x_locator1 ^ alpha420_2_x_locator2 ^ alpha420_3_x_locator3)), (~| (alpha419_0_x_locator0 ^ alpha419_1_x_locator1 ^ alpha419_2_x_locator2 ^ alpha419_3_x_locator3)), (~| (alpha418_0_x_locator0 ^ alpha418_1_x_locator1 ^ alpha418_2_x_locator2 ^ alpha418_3_x_locator3)), (~| (alpha417_0_x_locator0 ^ alpha417_1_x_locator1 ^ alpha417_2_x_locator2 ^ alpha417_3_x_locator3)), (~| (alpha416_0_x_locator0 ^ alpha416_1_x_locator1 ^ alpha416_2_x_locator2 ^ alpha416_3_x_locator3)), (~| (alpha415_0_x_locator0 ^ alpha415_1_x_locator1 ^ alpha415_2_x_locator2 ^ alpha415_3_x_locator3)), (~| (alpha414_0_x_locator0 ^ alpha414_1_x_locator1 ^ alpha414_2_x_locator2 ^ alpha414_3_x_locator3)), (~| (alpha413_0_x_locator0 ^ alpha413_1_x_locator1 ^ alpha413_2_x_locator2 ^ alpha413_3_x_locator3)), (~| (alpha412_0_x_locator0 ^ alpha412_1_x_locator1 ^ alpha412_2_x_locator2 ^ alpha412_3_x_locator3)), (~| (alpha411_0_x_locator0 ^ alpha411_1_x_locator1 ^ alpha411_2_x_locator2 ^ alpha411_3_x_locator3)), (~| (alpha410_0_x_locator0 ^ alpha410_1_x_locator1 ^ alpha410_2_x_locator2 ^ alpha410_3_x_locator3)), (~| (alpha409_0_x_locator0 ^ alpha409_1_x_locator1 ^ alpha409_2_x_locator2 ^ alpha409_3_x_locator3)), (~| (alpha408_0_x_locator0 ^ alpha408_1_x_locator1 ^ alpha408_2_x_locator2 ^ alpha408_3_x_locator3)), (~| (alpha407_0_x_locator0 ^ alpha407_1_x_locator1 ^ alpha407_2_x_locator2 ^ alpha407_3_x_locator3)), (~| (alpha406_0_x_locator0 ^ alpha406_1_x_locator1 ^ alpha406_2_x_locator2 ^ alpha406_3_x_locator3)), (~| (alpha405_0_x_locator0 ^ alpha405_1_x_locator1 ^ alpha405_2_x_locator2 ^ alpha405_3_x_locator3)), (~| (alpha404_0_x_locator0 ^ alpha404_1_x_locator1 ^ alpha404_2_x_locator2 ^ alpha404_3_x_locator3)), (~| (alpha403_0_x_locator0 ^ alpha403_1_x_locator1 ^ alpha403_2_x_locator2 ^ alpha403_3_x_locator3)), (~| (alpha402_0_x_locator0 ^ alpha402_1_x_locator1 ^ alpha402_2_x_locator2 ^ alpha402_3_x_locator3)), (~| (alpha401_0_x_locator0 ^ alpha401_1_x_locator1 ^ alpha401_2_x_locator2 ^ alpha401_3_x_locator3)), (~| (alpha400_0_x_locator0 ^ alpha400_1_x_locator1 ^ alpha400_2_x_locator2 ^ alpha400_3_x_locator3)), (~| (alpha399_0_x_locator0 ^ alpha399_1_x_locator1 ^ alpha399_2_x_locator2 ^ alpha399_3_x_locator3)), (~| (alpha398_0_x_locator0 ^ alpha398_1_x_locator1 ^ alpha398_2_x_locator2 ^ alpha398_3_x_locator3)), (~| (alpha397_0_x_locator0 ^ alpha397_1_x_locator1 ^ alpha397_2_x_locator2 ^ alpha397_3_x_locator3)), (~| (alpha396_0_x_locator0 ^ alpha396_1_x_locator1 ^ alpha396_2_x_locator2 ^ alpha396_3_x_locator3)), (~| (alpha395_0_x_locator0 ^ alpha395_1_x_locator1 ^ alpha395_2_x_locator2 ^ alpha395_3_x_locator3)), (~| (alpha394_0_x_locator0 ^ alpha394_1_x_locator1 ^ alpha394_2_x_locator2 ^ alpha394_3_x_locator3)), (~| (alpha393_0_x_locator0 ^ alpha393_1_x_locator1 ^ alpha393_2_x_locator2 ^ alpha393_3_x_locator3)), (~| (alpha392_0_x_locator0 ^ alpha392_1_x_locator1 ^ alpha392_2_x_locator2 ^ alpha392_3_x_locator3)), (~| (alpha391_0_x_locator0 ^ alpha391_1_x_locator1 ^ alpha391_2_x_locator2 ^ alpha391_3_x_locator3)), (~| (alpha390_0_x_locator0 ^ alpha390_1_x_locator1 ^ alpha390_2_x_locator2 ^ alpha390_3_x_locator3)), (~| (alpha389_0_x_locator0 ^ alpha389_1_x_locator1 ^ alpha389_2_x_locator2 ^ alpha389_3_x_locator3)), (~| (alpha388_0_x_locator0 ^ alpha388_1_x_locator1 ^ alpha388_2_x_locator2 ^ alpha388_3_x_locator3)), (~| (alpha387_0_x_locator0 ^ alpha387_1_x_locator1 ^ alpha387_2_x_locator2 ^ alpha387_3_x_locator3)), (~| (alpha386_0_x_locator0 ^ alpha386_1_x_locator1 ^ alpha386_2_x_locator2 ^ alpha386_3_x_locator3)), (~| (alpha385_0_x_locator0 ^ alpha385_1_x_locator1 ^ alpha385_2_x_locator2 ^ alpha385_3_x_locator3)), (~| (alpha384_0_x_locator0 ^ alpha384_1_x_locator1 ^ alpha384_2_x_locator2 ^ alpha384_3_x_locator3)), (~| (alpha383_0_x_locator0 ^ alpha383_1_x_locator1 ^ alpha383_2_x_locator2 ^ alpha383_3_x_locator3)), (~| (alpha382_0_x_locator0 ^ alpha382_1_x_locator1 ^ alpha382_2_x_locator2 ^ alpha382_3_x_locator3)), (~| (alpha381_0_x_locator0 ^ alpha381_1_x_locator1 ^ alpha381_2_x_locator2 ^ alpha381_3_x_locator3)), (~| (alpha380_0_x_locator0 ^ alpha380_1_x_locator1 ^ alpha380_2_x_locator2 ^ alpha380_3_x_locator3)), (~| (alpha379_0_x_locator0 ^ alpha379_1_x_locator1 ^ alpha379_2_x_locator2 ^ alpha379_3_x_locator3)), (~| (alpha378_0_x_locator0 ^ alpha378_1_x_locator1 ^ alpha378_2_x_locator2 ^ alpha378_3_x_locator3)), (~| (alpha377_0_x_locator0 ^ alpha377_1_x_locator1 ^ alpha377_2_x_locator2 ^ alpha377_3_x_locator3)), (~| (alpha376_0_x_locator0 ^ alpha376_1_x_locator1 ^ alpha376_2_x_locator2 ^ alpha376_3_x_locator3)), (~| (alpha375_0_x_locator0 ^ alpha375_1_x_locator1 ^ alpha375_2_x_locator2 ^ alpha375_3_x_locator3)), (~| (alpha374_0_x_locator0 ^ alpha374_1_x_locator1 ^ alpha374_2_x_locator2 ^ alpha374_3_x_locator3)), (~| (alpha373_0_x_locator0 ^ alpha373_1_x_locator1 ^ alpha373_2_x_locator2 ^ alpha373_3_x_locator3)), (~| (alpha372_0_x_locator0 ^ alpha372_1_x_locator1 ^ alpha372_2_x_locator2 ^ alpha372_3_x_locator3)), (~| (alpha371_0_x_locator0 ^ alpha371_1_x_locator1 ^ alpha371_2_x_locator2 ^ alpha371_3_x_locator3)), (~| (alpha370_0_x_locator0 ^ alpha370_1_x_locator1 ^ alpha370_2_x_locator2 ^ alpha370_3_x_locator3)), (~| (alpha369_0_x_locator0 ^ alpha369_1_x_locator1 ^ alpha369_2_x_locator2 ^ alpha369_3_x_locator3)), (~| (alpha368_0_x_locator0 ^ alpha368_1_x_locator1 ^ alpha368_2_x_locator2 ^ alpha368_3_x_locator3)), (~| (alpha367_0_x_locator0 ^ alpha367_1_x_locator1 ^ alpha367_2_x_locator2 ^ alpha367_3_x_locator3)), (~| (alpha366_0_x_locator0 ^ alpha366_1_x_locator1 ^ alpha366_2_x_locator2 ^ alpha366_3_x_locator3)), (~| (alpha365_0_x_locator0 ^ alpha365_1_x_locator1 ^ alpha365_2_x_locator2 ^ alpha365_3_x_locator3)), (~| (alpha364_0_x_locator0 ^ alpha364_1_x_locator1 ^ alpha364_2_x_locator2 ^ alpha364_3_x_locator3)), (~| (alpha363_0_x_locator0 ^ alpha363_1_x_locator1 ^ alpha363_2_x_locator2 ^ alpha363_3_x_locator3)), (~| (alpha362_0_x_locator0 ^ alpha362_1_x_locator1 ^ alpha362_2_x_locator2 ^ alpha362_3_x_locator3)), (~| (alpha361_0_x_locator0 ^ alpha361_1_x_locator1 ^ alpha361_2_x_locator2 ^ alpha361_3_x_locator3)), (~| (alpha360_0_x_locator0 ^ alpha360_1_x_locator1 ^ alpha360_2_x_locator2 ^ alpha360_3_x_locator3)), (~| (alpha359_0_x_locator0 ^ alpha359_1_x_locator1 ^ alpha359_2_x_locator2 ^ alpha359_3_x_locator3)), (~| (alpha358_0_x_locator0 ^ alpha358_1_x_locator1 ^ alpha358_2_x_locator2 ^ alpha358_3_x_locator3)), (~| (alpha357_0_x_locator0 ^ alpha357_1_x_locator1 ^ alpha357_2_x_locator2 ^ alpha357_3_x_locator3)), (~| (alpha356_0_x_locator0 ^ alpha356_1_x_locator1 ^ alpha356_2_x_locator2 ^ alpha356_3_x_locator3)), (~| (alpha355_0_x_locator0 ^ alpha355_1_x_locator1 ^ alpha355_2_x_locator2 ^ alpha355_3_x_locator3)), (~| (alpha354_0_x_locator0 ^ alpha354_1_x_locator1 ^ alpha354_2_x_locator2 ^ alpha354_3_x_locator3)), (~| (alpha353_0_x_locator0 ^ alpha353_1_x_locator1 ^ alpha353_2_x_locator2 ^ alpha353_3_x_locator3)), (~| (alpha352_0_x_locator0 ^ alpha352_1_x_locator1 ^ alpha352_2_x_locator2 ^ alpha352_3_x_locator3)), (~| (alpha351_0_x_locator0 ^ alpha351_1_x_locator1 ^ alpha351_2_x_locator2 ^ alpha351_3_x_locator3)), (~| (alpha350_0_x_locator0 ^ alpha350_1_x_locator1 ^ alpha350_2_x_locator2 ^ alpha350_3_x_locator3)), (~| (alpha349_0_x_locator0 ^ alpha349_1_x_locator1 ^ alpha349_2_x_locator2 ^ alpha349_3_x_locator3)), (~| (alpha348_0_x_locator0 ^ alpha348_1_x_locator1 ^ alpha348_2_x_locator2 ^ alpha348_3_x_locator3)), (~| (alpha347_0_x_locator0 ^ alpha347_1_x_locator1 ^ alpha347_2_x_locator2 ^ alpha347_3_x_locator3)), (~| (alpha346_0_x_locator0 ^ alpha346_1_x_locator1 ^ alpha346_2_x_locator2 ^ alpha346_3_x_locator3)), (~| (alpha345_0_x_locator0 ^ alpha345_1_x_locator1 ^ alpha345_2_x_locator2 ^ alpha345_3_x_locator3)), (~| (alpha344_0_x_locator0 ^ alpha344_1_x_locator1 ^ alpha344_2_x_locator2 ^ alpha344_3_x_locator3)), (~| (alpha343_0_x_locator0 ^ alpha343_1_x_locator1 ^ alpha343_2_x_locator2 ^ alpha343_3_x_locator3)), (~| (alpha342_0_x_locator0 ^ alpha342_1_x_locator1 ^ alpha342_2_x_locator2 ^ alpha342_3_x_locator3)), (~| (alpha341_0_x_locator0 ^ alpha341_1_x_locator1 ^ alpha341_2_x_locator2 ^ alpha341_3_x_locator3)), (~| (alpha340_0_x_locator0 ^ alpha340_1_x_locator1 ^ alpha340_2_x_locator2 ^ alpha340_3_x_locator3)), (~| (alpha339_0_x_locator0 ^ alpha339_1_x_locator1 ^ alpha339_2_x_locator2 ^ alpha339_3_x_locator3)), (~| (alpha338_0_x_locator0 ^ alpha338_1_x_locator1 ^ alpha338_2_x_locator2 ^ alpha338_3_x_locator3)), (~| (alpha337_0_x_locator0 ^ alpha337_1_x_locator1 ^ alpha337_2_x_locator2 ^ alpha337_3_x_locator3)), (~| (alpha336_0_x_locator0 ^ alpha336_1_x_locator1 ^ alpha336_2_x_locator2 ^ alpha336_3_x_locator3)), (~| (alpha335_0_x_locator0 ^ alpha335_1_x_locator1 ^ alpha335_2_x_locator2 ^ alpha335_3_x_locator3)), (~| (alpha334_0_x_locator0 ^ alpha334_1_x_locator1 ^ alpha334_2_x_locator2 ^ alpha334_3_x_locator3)), (~| (alpha333_0_x_locator0 ^ alpha333_1_x_locator1 ^ alpha333_2_x_locator2 ^ alpha333_3_x_locator3)), (~| (alpha332_0_x_locator0 ^ alpha332_1_x_locator1 ^ alpha332_2_x_locator2 ^ alpha332_3_x_locator3)), (~| (alpha331_0_x_locator0 ^ alpha331_1_x_locator1 ^ alpha331_2_x_locator2 ^ alpha331_3_x_locator3)), (~| (alpha330_0_x_locator0 ^ alpha330_1_x_locator1 ^ alpha330_2_x_locator2 ^ alpha330_3_x_locator3)), (~| (alpha329_0_x_locator0 ^ alpha329_1_x_locator1 ^ alpha329_2_x_locator2 ^ alpha329_3_x_locator3)), (~| (alpha328_0_x_locator0 ^ alpha328_1_x_locator1 ^ alpha328_2_x_locator2 ^ alpha328_3_x_locator3)), (~| (alpha327_0_x_locator0 ^ alpha327_1_x_locator1 ^ alpha327_2_x_locator2 ^ alpha327_3_x_locator3)), (~| (alpha326_0_x_locator0 ^ alpha326_1_x_locator1 ^ alpha326_2_x_locator2 ^ alpha326_3_x_locator3)), (~| (alpha325_0_x_locator0 ^ alpha325_1_x_locator1 ^ alpha325_2_x_locator2 ^ alpha325_3_x_locator3)), (~| (alpha324_0_x_locator0 ^ alpha324_1_x_locator1 ^ alpha324_2_x_locator2 ^ alpha324_3_x_locator3)), (~| (alpha323_0_x_locator0 ^ alpha323_1_x_locator1 ^ alpha323_2_x_locator2 ^ alpha323_3_x_locator3)), (~| (alpha322_0_x_locator0 ^ alpha322_1_x_locator1 ^ alpha322_2_x_locator2 ^ alpha322_3_x_locator3)), (~| (alpha321_0_x_locator0 ^ alpha321_1_x_locator1 ^ alpha321_2_x_locator2 ^ alpha321_3_x_locator3)), (~| (alpha320_0_x_locator0 ^ alpha320_1_x_locator1 ^ alpha320_2_x_locator2 ^ alpha320_3_x_locator3)), (~| (alpha319_0_x_locator0 ^ alpha319_1_x_locator1 ^ alpha319_2_x_locator2 ^ alpha319_3_x_locator3)), (~| (alpha318_0_x_locator0 ^ alpha318_1_x_locator1 ^ alpha318_2_x_locator2 ^ alpha318_3_x_locator3)), (~| (alpha317_0_x_locator0 ^ alpha317_1_x_locator1 ^ alpha317_2_x_locator2 ^ alpha317_3_x_locator3)), (~| (alpha316_0_x_locator0 ^ alpha316_1_x_locator1 ^ alpha316_2_x_locator2 ^ alpha316_3_x_locator3)), (~| (alpha315_0_x_locator0 ^ alpha315_1_x_locator1 ^ alpha315_2_x_locator2 ^ alpha315_3_x_locator3)), (~| (alpha314_0_x_locator0 ^ alpha314_1_x_locator1 ^ alpha314_2_x_locator2 ^ alpha314_3_x_locator3)), (~| (alpha313_0_x_locator0 ^ alpha313_1_x_locator1 ^ alpha313_2_x_locator2 ^ alpha313_3_x_locator3)), (~| (alpha312_0_x_locator0 ^ alpha312_1_x_locator1 ^ alpha312_2_x_locator2 ^ alpha312_3_x_locator3)), (~| (alpha311_0_x_locator0 ^ alpha311_1_x_locator1 ^ alpha311_2_x_locator2 ^ alpha311_3_x_locator3)), (~| (alpha310_0_x_locator0 ^ alpha310_1_x_locator1 ^ alpha310_2_x_locator2 ^ alpha310_3_x_locator3)), (~| (alpha309_0_x_locator0 ^ alpha309_1_x_locator1 ^ alpha309_2_x_locator2 ^ alpha309_3_x_locator3)), (~| (alpha308_0_x_locator0 ^ alpha308_1_x_locator1 ^ alpha308_2_x_locator2 ^ alpha308_3_x_locator3)), (~| (alpha307_0_x_locator0 ^ alpha307_1_x_locator1 ^ alpha307_2_x_locator2 ^ alpha307_3_x_locator3)), (~| (alpha306_0_x_locator0 ^ alpha306_1_x_locator1 ^ alpha306_2_x_locator2 ^ alpha306_3_x_locator3)), (~| (alpha305_0_x_locator0 ^ alpha305_1_x_locator1 ^ alpha305_2_x_locator2 ^ alpha305_3_x_locator3)), (~| (alpha304_0_x_locator0 ^ alpha304_1_x_locator1 ^ alpha304_2_x_locator2 ^ alpha304_3_x_locator3)), (~| (alpha303_0_x_locator0 ^ alpha303_1_x_locator1 ^ alpha303_2_x_locator2 ^ alpha303_3_x_locator3)), (~| (alpha302_0_x_locator0 ^ alpha302_1_x_locator1 ^ alpha302_2_x_locator2 ^ alpha302_3_x_locator3)), (~| (alpha301_0_x_locator0 ^ alpha301_1_x_locator1 ^ alpha301_2_x_locator2 ^ alpha301_3_x_locator3)), (~| (alpha300_0_x_locator0 ^ alpha300_1_x_locator1 ^ alpha300_2_x_locator2 ^ alpha300_3_x_locator3)), (~| (alpha299_0_x_locator0 ^ alpha299_1_x_locator1 ^ alpha299_2_x_locator2 ^ alpha299_3_x_locator3)), (~| (alpha298_0_x_locator0 ^ alpha298_1_x_locator1 ^ alpha298_2_x_locator2 ^ alpha298_3_x_locator3)), (~| (alpha297_0_x_locator0 ^ alpha297_1_x_locator1 ^ alpha297_2_x_locator2 ^ alpha297_3_x_locator3)), (~| (alpha296_0_x_locator0 ^ alpha296_1_x_locator1 ^ alpha296_2_x_locator2 ^ alpha296_3_x_locator3)), (~| (alpha295_0_x_locator0 ^ alpha295_1_x_locator1 ^ alpha295_2_x_locator2 ^ alpha295_3_x_locator3)), (~| (alpha294_0_x_locator0 ^ alpha294_1_x_locator1 ^ alpha294_2_x_locator2 ^ alpha294_3_x_locator3)), (~| (alpha293_0_x_locator0 ^ alpha293_1_x_locator1 ^ alpha293_2_x_locator2 ^ alpha293_3_x_locator3)), (~| (alpha292_0_x_locator0 ^ alpha292_1_x_locator1 ^ alpha292_2_x_locator2 ^ alpha292_3_x_locator3)), (~| (alpha291_0_x_locator0 ^ alpha291_1_x_locator1 ^ alpha291_2_x_locator2 ^ alpha291_3_x_locator3)), (~| (alpha290_0_x_locator0 ^ alpha290_1_x_locator1 ^ alpha290_2_x_locator2 ^ alpha290_3_x_locator3)), (~| (alpha289_0_x_locator0 ^ alpha289_1_x_locator1 ^ alpha289_2_x_locator2 ^ alpha289_3_x_locator3)), (~| (alpha288_0_x_locator0 ^ alpha288_1_x_locator1 ^ alpha288_2_x_locator2 ^ alpha288_3_x_locator3)), (~| (alpha287_0_x_locator0 ^ alpha287_1_x_locator1 ^ alpha287_2_x_locator2 ^ alpha287_3_x_locator3)), (~| (alpha286_0_x_locator0 ^ alpha286_1_x_locator1 ^ alpha286_2_x_locator2 ^ alpha286_3_x_locator3)), (~| (alpha285_0_x_locator0 ^ alpha285_1_x_locator1 ^ alpha285_2_x_locator2 ^ alpha285_3_x_locator3)), (~| (alpha284_0_x_locator0 ^ alpha284_1_x_locator1 ^ alpha284_2_x_locator2 ^ alpha284_3_x_locator3)), (~| (alpha283_0_x_locator0 ^ alpha283_1_x_locator1 ^ alpha283_2_x_locator2 ^ alpha283_3_x_locator3)), (~| (alpha282_0_x_locator0 ^ alpha282_1_x_locator1 ^ alpha282_2_x_locator2 ^ alpha282_3_x_locator3)), (~| (alpha281_0_x_locator0 ^ alpha281_1_x_locator1 ^ alpha281_2_x_locator2 ^ alpha281_3_x_locator3)), (~| (alpha280_0_x_locator0 ^ alpha280_1_x_locator1 ^ alpha280_2_x_locator2 ^ alpha280_3_x_locator3)), (~| (alpha279_0_x_locator0 ^ alpha279_1_x_locator1 ^ alpha279_2_x_locator2 ^ alpha279_3_x_locator3)), (~| (alpha278_0_x_locator0 ^ alpha278_1_x_locator1 ^ alpha278_2_x_locator2 ^ alpha278_3_x_locator3)), (~| (alpha277_0_x_locator0 ^ alpha277_1_x_locator1 ^ alpha277_2_x_locator2 ^ alpha277_3_x_locator3)), (~| (alpha276_0_x_locator0 ^ alpha276_1_x_locator1 ^ alpha276_2_x_locator2 ^ alpha276_3_x_locator3)), (~| (alpha275_0_x_locator0 ^ alpha275_1_x_locator1 ^ alpha275_2_x_locator2 ^ alpha275_3_x_locator3)), (~| (alpha274_0_x_locator0 ^ alpha274_1_x_locator1 ^ alpha274_2_x_locator2 ^ alpha274_3_x_locator3)), (~| (alpha273_0_x_locator0 ^ alpha273_1_x_locator1 ^ alpha273_2_x_locator2 ^ alpha273_3_x_locator3)), (~| (alpha272_0_x_locator0 ^ alpha272_1_x_locator1 ^ alpha272_2_x_locator2 ^ alpha272_3_x_locator3)), (~| (alpha271_0_x_locator0 ^ alpha271_1_x_locator1 ^ alpha271_2_x_locator2 ^ alpha271_3_x_locator3)), (~| (alpha270_0_x_locator0 ^ alpha270_1_x_locator1 ^ alpha270_2_x_locator2 ^ alpha270_3_x_locator3)), (~| (alpha269_0_x_locator0 ^ alpha269_1_x_locator1 ^ alpha269_2_x_locator2 ^ alpha269_3_x_locator3)), (~| (alpha268_0_x_locator0 ^ alpha268_1_x_locator1 ^ alpha268_2_x_locator2 ^ alpha268_3_x_locator3)), (~| (alpha267_0_x_locator0 ^ alpha267_1_x_locator1 ^ alpha267_2_x_locator2 ^ alpha267_3_x_locator3)), (~| (alpha266_0_x_locator0 ^ alpha266_1_x_locator1 ^ alpha266_2_x_locator2 ^ alpha266_3_x_locator3)), (~| (alpha265_0_x_locator0 ^ alpha265_1_x_locator1 ^ alpha265_2_x_locator2 ^ alpha265_3_x_locator3)), (~| (alpha264_0_x_locator0 ^ alpha264_1_x_locator1 ^ alpha264_2_x_locator2 ^ alpha264_3_x_locator3)), (~| (alpha263_0_x_locator0 ^ alpha263_1_x_locator1 ^ alpha263_2_x_locator2 ^ alpha263_3_x_locator3)), (~| (alpha262_0_x_locator0 ^ alpha262_1_x_locator1 ^ alpha262_2_x_locator2 ^ alpha262_3_x_locator3)), (~| (alpha261_0_x_locator0 ^ alpha261_1_x_locator1 ^ alpha261_2_x_locator2 ^ alpha261_3_x_locator3)), (~| (alpha260_0_x_locator0 ^ alpha260_1_x_locator1 ^ alpha260_2_x_locator2 ^ alpha260_3_x_locator3)), (~| (alpha259_0_x_locator0 ^ alpha259_1_x_locator1 ^ alpha259_2_x_locator2 ^ alpha259_3_x_locator3)), (~| (alpha258_0_x_locator0 ^ alpha258_1_x_locator1 ^ alpha258_2_x_locator2 ^ alpha258_3_x_locator3)), (~| (alpha257_0_x_locator0 ^ alpha257_1_x_locator1 ^ alpha257_2_x_locator2 ^ alpha257_3_x_locator3)), (~| (alpha256_0_x_locator0 ^ alpha256_1_x_locator1 ^ alpha256_2_x_locator2 ^ alpha256_3_x_locator3)), (~| (alpha255_0_x_locator0 ^ alpha255_1_x_locator1 ^ alpha255_2_x_locator2 ^ alpha255_3_x_locator3)), (~| (alpha254_0_x_locator0 ^ alpha254_1_x_locator1 ^ alpha254_2_x_locator2 ^ alpha254_3_x_locator3)), (~| (alpha253_0_x_locator0 ^ alpha253_1_x_locator1 ^ alpha253_2_x_locator2 ^ alpha253_3_x_locator3)), (~| (alpha252_0_x_locator0 ^ alpha252_1_x_locator1 ^ alpha252_2_x_locator2 ^ alpha252_3_x_locator3)), (~| (alpha251_0_x_locator0 ^ alpha251_1_x_locator1 ^ alpha251_2_x_locator2 ^ alpha251_3_x_locator3)), (~| (alpha250_0_x_locator0 ^ alpha250_1_x_locator1 ^ alpha250_2_x_locator2 ^ alpha250_3_x_locator3)), (~| (alpha249_0_x_locator0 ^ alpha249_1_x_locator1 ^ alpha249_2_x_locator2 ^ alpha249_3_x_locator3)), (~| (alpha248_0_x_locator0 ^ alpha248_1_x_locator1 ^ alpha248_2_x_locator2 ^ alpha248_3_x_locator3)), (~| (alpha247_0_x_locator0 ^ alpha247_1_x_locator1 ^ alpha247_2_x_locator2 ^ alpha247_3_x_locator3)), (~| (alpha246_0_x_locator0 ^ alpha246_1_x_locator1 ^ alpha246_2_x_locator2 ^ alpha246_3_x_locator3)), (~| (alpha245_0_x_locator0 ^ alpha245_1_x_locator1 ^ alpha245_2_x_locator2 ^ alpha245_3_x_locator3)), (~| (alpha244_0_x_locator0 ^ alpha244_1_x_locator1 ^ alpha244_2_x_locator2 ^ alpha244_3_x_locator3)), (~| (alpha243_0_x_locator0 ^ alpha243_1_x_locator1 ^ alpha243_2_x_locator2 ^ alpha243_3_x_locator3)), (~| (alpha242_0_x_locator0 ^ alpha242_1_x_locator1 ^ alpha242_2_x_locator2 ^ alpha242_3_x_locator3)), (~| (alpha241_0_x_locator0 ^ alpha241_1_x_locator1 ^ alpha241_2_x_locator2 ^ alpha241_3_x_locator3)), (~| (alpha240_0_x_locator0 ^ alpha240_1_x_locator1 ^ alpha240_2_x_locator2 ^ alpha240_3_x_locator3)), (~| (alpha239_0_x_locator0 ^ alpha239_1_x_locator1 ^ alpha239_2_x_locator2 ^ alpha239_3_x_locator3)), (~| (alpha238_0_x_locator0 ^ alpha238_1_x_locator1 ^ alpha238_2_x_locator2 ^ alpha238_3_x_locator3)), (~| (alpha237_0_x_locator0 ^ alpha237_1_x_locator1 ^ alpha237_2_x_locator2 ^ alpha237_3_x_locator3)), (~| (alpha236_0_x_locator0 ^ alpha236_1_x_locator1 ^ alpha236_2_x_locator2 ^ alpha236_3_x_locator3)), (~| (alpha235_0_x_locator0 ^ alpha235_1_x_locator1 ^ alpha235_2_x_locator2 ^ alpha235_3_x_locator3)), (~| (alpha234_0_x_locator0 ^ alpha234_1_x_locator1 ^ alpha234_2_x_locator2 ^ alpha234_3_x_locator3)), (~| (alpha233_0_x_locator0 ^ alpha233_1_x_locator1 ^ alpha233_2_x_locator2 ^ alpha233_3_x_locator3)), (~| (alpha232_0_x_locator0 ^ alpha232_1_x_locator1 ^ alpha232_2_x_locator2 ^ alpha232_3_x_locator3)), (~| (alpha231_0_x_locator0 ^ alpha231_1_x_locator1 ^ alpha231_2_x_locator2 ^ alpha231_3_x_locator3)), (~| (alpha230_0_x_locator0 ^ alpha230_1_x_locator1 ^ alpha230_2_x_locator2 ^ alpha230_3_x_locator3)), (~| (alpha229_0_x_locator0 ^ alpha229_1_x_locator1 ^ alpha229_2_x_locator2 ^ alpha229_3_x_locator3)), (~| (alpha228_0_x_locator0 ^ alpha228_1_x_locator1 ^ alpha228_2_x_locator2 ^ alpha228_3_x_locator3)), (~| (alpha227_0_x_locator0 ^ alpha227_1_x_locator1 ^ alpha227_2_x_locator2 ^ alpha227_3_x_locator3)), (~| (alpha226_0_x_locator0 ^ alpha226_1_x_locator1 ^ alpha226_2_x_locator2 ^ alpha226_3_x_locator3)), (~| (alpha225_0_x_locator0 ^ alpha225_1_x_locator1 ^ alpha225_2_x_locator2 ^ alpha225_3_x_locator3)), (~| (alpha224_0_x_locator0 ^ alpha224_1_x_locator1 ^ alpha224_2_x_locator2 ^ alpha224_3_x_locator3)), (~| (alpha223_0_x_locator0 ^ alpha223_1_x_locator1 ^ alpha223_2_x_locator2 ^ alpha223_3_x_locator3)), (~| (alpha222_0_x_locator0 ^ alpha222_1_x_locator1 ^ alpha222_2_x_locator2 ^ alpha222_3_x_locator3)), (~| (alpha221_0_x_locator0 ^ alpha221_1_x_locator1 ^ alpha221_2_x_locator2 ^ alpha221_3_x_locator3)), (~| (alpha220_0_x_locator0 ^ alpha220_1_x_locator1 ^ alpha220_2_x_locator2 ^ alpha220_3_x_locator3)), (~| (alpha219_0_x_locator0 ^ alpha219_1_x_locator1 ^ alpha219_2_x_locator2 ^ alpha219_3_x_locator3)), (~| (alpha218_0_x_locator0 ^ alpha218_1_x_locator1 ^ alpha218_2_x_locator2 ^ alpha218_3_x_locator3)), (~| (alpha217_0_x_locator0 ^ alpha217_1_x_locator1 ^ alpha217_2_x_locator2 ^ alpha217_3_x_locator3)), (~| (alpha216_0_x_locator0 ^ alpha216_1_x_locator1 ^ alpha216_2_x_locator2 ^ alpha216_3_x_locator3)), (~| (alpha215_0_x_locator0 ^ alpha215_1_x_locator1 ^ alpha215_2_x_locator2 ^ alpha215_3_x_locator3)), (~| (alpha214_0_x_locator0 ^ alpha214_1_x_locator1 ^ alpha214_2_x_locator2 ^ alpha214_3_x_locator3)), (~| (alpha213_0_x_locator0 ^ alpha213_1_x_locator1 ^ alpha213_2_x_locator2 ^ alpha213_3_x_locator3)), (~| (alpha212_0_x_locator0 ^ alpha212_1_x_locator1 ^ alpha212_2_x_locator2 ^ alpha212_3_x_locator3)), (~| (alpha211_0_x_locator0 ^ alpha211_1_x_locator1 ^ alpha211_2_x_locator2 ^ alpha211_3_x_locator3)), (~| (alpha210_0_x_locator0 ^ alpha210_1_x_locator1 ^ alpha210_2_x_locator2 ^ alpha210_3_x_locator3)), (~| (alpha209_0_x_locator0 ^ alpha209_1_x_locator1 ^ alpha209_2_x_locator2 ^ alpha209_3_x_locator3)), (~| (alpha208_0_x_locator0 ^ alpha208_1_x_locator1 ^ alpha208_2_x_locator2 ^ alpha208_3_x_locator3)), (~| (alpha207_0_x_locator0 ^ alpha207_1_x_locator1 ^ alpha207_2_x_locator2 ^ alpha207_3_x_locator3)), (~| (alpha206_0_x_locator0 ^ alpha206_1_x_locator1 ^ alpha206_2_x_locator2 ^ alpha206_3_x_locator3)), (~| (alpha205_0_x_locator0 ^ alpha205_1_x_locator1 ^ alpha205_2_x_locator2 ^ alpha205_3_x_locator3)), (~| (alpha204_0_x_locator0 ^ alpha204_1_x_locator1 ^ alpha204_2_x_locator2 ^ alpha204_3_x_locator3)), (~| (alpha203_0_x_locator0 ^ alpha203_1_x_locator1 ^ alpha203_2_x_locator2 ^ alpha203_3_x_locator3)), (~| (alpha202_0_x_locator0 ^ alpha202_1_x_locator1 ^ alpha202_2_x_locator2 ^ alpha202_3_x_locator3)), (~| (alpha201_0_x_locator0 ^ alpha201_1_x_locator1 ^ alpha201_2_x_locator2 ^ alpha201_3_x_locator3)), (~| (alpha200_0_x_locator0 ^ alpha200_1_x_locator1 ^ alpha200_2_x_locator2 ^ alpha200_3_x_locator3)), (~| (alpha199_0_x_locator0 ^ alpha199_1_x_locator1 ^ alpha199_2_x_locator2 ^ alpha199_3_x_locator3)), (~| (alpha198_0_x_locator0 ^ alpha198_1_x_locator1 ^ alpha198_2_x_locator2 ^ alpha198_3_x_locator3)), (~| (alpha197_0_x_locator0 ^ alpha197_1_x_locator1 ^ alpha197_2_x_locator2 ^ alpha197_3_x_locator3)), (~| (alpha196_0_x_locator0 ^ alpha196_1_x_locator1 ^ alpha196_2_x_locator2 ^ alpha196_3_x_locator3)), (~| (alpha195_0_x_locator0 ^ alpha195_1_x_locator1 ^ alpha195_2_x_locator2 ^ alpha195_3_x_locator3)), (~| (alpha194_0_x_locator0 ^ alpha194_1_x_locator1 ^ alpha194_2_x_locator2 ^ alpha194_3_x_locator3)), (~| (alpha193_0_x_locator0 ^ alpha193_1_x_locator1 ^ alpha193_2_x_locator2 ^ alpha193_3_x_locator3)), (~| (alpha192_0_x_locator0 ^ alpha192_1_x_locator1 ^ alpha192_2_x_locator2 ^ alpha192_3_x_locator3)), (~| (alpha191_0_x_locator0 ^ alpha191_1_x_locator1 ^ alpha191_2_x_locator2 ^ alpha191_3_x_locator3)), (~| (alpha190_0_x_locator0 ^ alpha190_1_x_locator1 ^ alpha190_2_x_locator2 ^ alpha190_3_x_locator3)), (~| (alpha189_0_x_locator0 ^ alpha189_1_x_locator1 ^ alpha189_2_x_locator2 ^ alpha189_3_x_locator3)), (~| (alpha188_0_x_locator0 ^ alpha188_1_x_locator1 ^ alpha188_2_x_locator2 ^ alpha188_3_x_locator3)), (~| (alpha187_0_x_locator0 ^ alpha187_1_x_locator1 ^ alpha187_2_x_locator2 ^ alpha187_3_x_locator3)), (~| (alpha186_0_x_locator0 ^ alpha186_1_x_locator1 ^ alpha186_2_x_locator2 ^ alpha186_3_x_locator3)), (~| (alpha185_0_x_locator0 ^ alpha185_1_x_locator1 ^ alpha185_2_x_locator2 ^ alpha185_3_x_locator3)), (~| (alpha184_0_x_locator0 ^ alpha184_1_x_locator1 ^ alpha184_2_x_locator2 ^ alpha184_3_x_locator3)), (~| (alpha183_0_x_locator0 ^ alpha183_1_x_locator1 ^ alpha183_2_x_locator2 ^ alpha183_3_x_locator3)), (~| (alpha182_0_x_locator0 ^ alpha182_1_x_locator1 ^ alpha182_2_x_locator2 ^ alpha182_3_x_locator3)), (~| (alpha181_0_x_locator0 ^ alpha181_1_x_locator1 ^ alpha181_2_x_locator2 ^ alpha181_3_x_locator3)), (~| (alpha180_0_x_locator0 ^ alpha180_1_x_locator1 ^ alpha180_2_x_locator2 ^ alpha180_3_x_locator3)), (~| (alpha179_0_x_locator0 ^ alpha179_1_x_locator1 ^ alpha179_2_x_locator2 ^ alpha179_3_x_locator3)), (~| (alpha178_0_x_locator0 ^ alpha178_1_x_locator1 ^ alpha178_2_x_locator2 ^ alpha178_3_x_locator3)), (~| (alpha177_0_x_locator0 ^ alpha177_1_x_locator1 ^ alpha177_2_x_locator2 ^ alpha177_3_x_locator3)), (~| (alpha176_0_x_locator0 ^ alpha176_1_x_locator1 ^ alpha176_2_x_locator2 ^ alpha176_3_x_locator3)), (~| (alpha175_0_x_locator0 ^ alpha175_1_x_locator1 ^ alpha175_2_x_locator2 ^ alpha175_3_x_locator3)), (~| (alpha174_0_x_locator0 ^ alpha174_1_x_locator1 ^ alpha174_2_x_locator2 ^ alpha174_3_x_locator3)), (~| (alpha173_0_x_locator0 ^ alpha173_1_x_locator1 ^ alpha173_2_x_locator2 ^ alpha173_3_x_locator3)), (~| (alpha172_0_x_locator0 ^ alpha172_1_x_locator1 ^ alpha172_2_x_locator2 ^ alpha172_3_x_locator3)), (~| (alpha171_0_x_locator0 ^ alpha171_1_x_locator1 ^ alpha171_2_x_locator2 ^ alpha171_3_x_locator3)), (~| (alpha170_0_x_locator0 ^ alpha170_1_x_locator1 ^ alpha170_2_x_locator2 ^ alpha170_3_x_locator3)), (~| (alpha169_0_x_locator0 ^ alpha169_1_x_locator1 ^ alpha169_2_x_locator2 ^ alpha169_3_x_locator3)), (~| (alpha168_0_x_locator0 ^ alpha168_1_x_locator1 ^ alpha168_2_x_locator2 ^ alpha168_3_x_locator3)), (~| (alpha167_0_x_locator0 ^ alpha167_1_x_locator1 ^ alpha167_2_x_locator2 ^ alpha167_3_x_locator3)), (~| (alpha166_0_x_locator0 ^ alpha166_1_x_locator1 ^ alpha166_2_x_locator2 ^ alpha166_3_x_locator3)), (~| (alpha165_0_x_locator0 ^ alpha165_1_x_locator1 ^ alpha165_2_x_locator2 ^ alpha165_3_x_locator3)), (~| (alpha164_0_x_locator0 ^ alpha164_1_x_locator1 ^ alpha164_2_x_locator2 ^ alpha164_3_x_locator3)), (~| (alpha163_0_x_locator0 ^ alpha163_1_x_locator1 ^ alpha163_2_x_locator2 ^ alpha163_3_x_locator3)), (~| (alpha162_0_x_locator0 ^ alpha162_1_x_locator1 ^ alpha162_2_x_locator2 ^ alpha162_3_x_locator3)), (~| (alpha161_0_x_locator0 ^ alpha161_1_x_locator1 ^ alpha161_2_x_locator2 ^ alpha161_3_x_locator3)), (~| (alpha160_0_x_locator0 ^ alpha160_1_x_locator1 ^ alpha160_2_x_locator2 ^ alpha160_3_x_locator3)), (~| (alpha159_0_x_locator0 ^ alpha159_1_x_locator1 ^ alpha159_2_x_locator2 ^ alpha159_3_x_locator3)), (~| (alpha158_0_x_locator0 ^ alpha158_1_x_locator1 ^ alpha158_2_x_locator2 ^ alpha158_3_x_locator3)), (~| (alpha157_0_x_locator0 ^ alpha157_1_x_locator1 ^ alpha157_2_x_locator2 ^ alpha157_3_x_locator3)), (~| (alpha156_0_x_locator0 ^ alpha156_1_x_locator1 ^ alpha156_2_x_locator2 ^ alpha156_3_x_locator3)), (~| (alpha155_0_x_locator0 ^ alpha155_1_x_locator1 ^ alpha155_2_x_locator2 ^ alpha155_3_x_locator3)), (~| (alpha154_0_x_locator0 ^ alpha154_1_x_locator1 ^ alpha154_2_x_locator2 ^ alpha154_3_x_locator3)), (~| (alpha153_0_x_locator0 ^ alpha153_1_x_locator1 ^ alpha153_2_x_locator2 ^ alpha153_3_x_locator3)), (~| (alpha152_0_x_locator0 ^ alpha152_1_x_locator1 ^ alpha152_2_x_locator2 ^ alpha152_3_x_locator3)), (~| (alpha151_0_x_locator0 ^ alpha151_1_x_locator1 ^ alpha151_2_x_locator2 ^ alpha151_3_x_locator3)), (~| (alpha150_0_x_locator0 ^ alpha150_1_x_locator1 ^ alpha150_2_x_locator2 ^ alpha150_3_x_locator3)), (~| (alpha149_0_x_locator0 ^ alpha149_1_x_locator1 ^ alpha149_2_x_locator2 ^ alpha149_3_x_locator3)), (~| (alpha148_0_x_locator0 ^ alpha148_1_x_locator1 ^ alpha148_2_x_locator2 ^ alpha148_3_x_locator3)), (~| (alpha147_0_x_locator0 ^ alpha147_1_x_locator1 ^ alpha147_2_x_locator2 ^ alpha147_3_x_locator3)), (~| (alpha146_0_x_locator0 ^ alpha146_1_x_locator1 ^ alpha146_2_x_locator2 ^ alpha146_3_x_locator3)), (~| (alpha145_0_x_locator0 ^ alpha145_1_x_locator1 ^ alpha145_2_x_locator2 ^ alpha145_3_x_locator3)), (~| (alpha144_0_x_locator0 ^ alpha144_1_x_locator1 ^ alpha144_2_x_locator2 ^ alpha144_3_x_locator3)), (~| (alpha143_0_x_locator0 ^ alpha143_1_x_locator1 ^ alpha143_2_x_locator2 ^ alpha143_3_x_locator3)), (~| (alpha142_0_x_locator0 ^ alpha142_1_x_locator1 ^ alpha142_2_x_locator2 ^ alpha142_3_x_locator3)), (~| (alpha141_0_x_locator0 ^ alpha141_1_x_locator1 ^ alpha141_2_x_locator2 ^ alpha141_3_x_locator3)), (~| (alpha140_0_x_locator0 ^ alpha140_1_x_locator1 ^ alpha140_2_x_locator2 ^ alpha140_3_x_locator3)), (~| (alpha139_0_x_locator0 ^ alpha139_1_x_locator1 ^ alpha139_2_x_locator2 ^ alpha139_3_x_locator3)), (~| (alpha138_0_x_locator0 ^ alpha138_1_x_locator1 ^ alpha138_2_x_locator2 ^ alpha138_3_x_locator3)), (~| (alpha137_0_x_locator0 ^ alpha137_1_x_locator1 ^ alpha137_2_x_locator2 ^ alpha137_3_x_locator3)), (~| (alpha136_0_x_locator0 ^ alpha136_1_x_locator1 ^ alpha136_2_x_locator2 ^ alpha136_3_x_locator3)), (~| (alpha135_0_x_locator0 ^ alpha135_1_x_locator1 ^ alpha135_2_x_locator2 ^ alpha135_3_x_locator3)), (~| (alpha134_0_x_locator0 ^ alpha134_1_x_locator1 ^ alpha134_2_x_locator2 ^ alpha134_3_x_locator3)), (~| (alpha133_0_x_locator0 ^ alpha133_1_x_locator1 ^ alpha133_2_x_locator2 ^ alpha133_3_x_locator3)), (~| (alpha132_0_x_locator0 ^ alpha132_1_x_locator1 ^ alpha132_2_x_locator2 ^ alpha132_3_x_locator3)), (~| (alpha131_0_x_locator0 ^ alpha131_1_x_locator1 ^ alpha131_2_x_locator2 ^ alpha131_3_x_locator3)), (~| (alpha130_0_x_locator0 ^ alpha130_1_x_locator1 ^ alpha130_2_x_locator2 ^ alpha130_3_x_locator3)), (~| (alpha129_0_x_locator0 ^ alpha129_1_x_locator1 ^ alpha129_2_x_locator2 ^ alpha129_3_x_locator3)), (~| (alpha128_0_x_locator0 ^ alpha128_1_x_locator1 ^ alpha128_2_x_locator2 ^ alpha128_3_x_locator3)), (~| (alpha127_0_x_locator0 ^ alpha127_1_x_locator1 ^ alpha127_2_x_locator2 ^ alpha127_3_x_locator3)), (~| (alpha126_0_x_locator0 ^ alpha126_1_x_locator1 ^ alpha126_2_x_locator2 ^ alpha126_3_x_locator3)), (~| (alpha125_0_x_locator0 ^ alpha125_1_x_locator1 ^ alpha125_2_x_locator2 ^ alpha125_3_x_locator3)), (~| (alpha124_0_x_locator0 ^ alpha124_1_x_locator1 ^ alpha124_2_x_locator2 ^ alpha124_3_x_locator3)), (~| (alpha123_0_x_locator0 ^ alpha123_1_x_locator1 ^ alpha123_2_x_locator2 ^ alpha123_3_x_locator3)), (~| (alpha122_0_x_locator0 ^ alpha122_1_x_locator1 ^ alpha122_2_x_locator2 ^ alpha122_3_x_locator3)), (~| (alpha121_0_x_locator0 ^ alpha121_1_x_locator1 ^ alpha121_2_x_locator2 ^ alpha121_3_x_locator3)), (~| (alpha120_0_x_locator0 ^ alpha120_1_x_locator1 ^ alpha120_2_x_locator2 ^ alpha120_3_x_locator3)), (~| (alpha119_0_x_locator0 ^ alpha119_1_x_locator1 ^ alpha119_2_x_locator2 ^ alpha119_3_x_locator3)), (~| (alpha118_0_x_locator0 ^ alpha118_1_x_locator1 ^ alpha118_2_x_locator2 ^ alpha118_3_x_locator3)), (~| (alpha117_0_x_locator0 ^ alpha117_1_x_locator1 ^ alpha117_2_x_locator2 ^ alpha117_3_x_locator3)), (~| (alpha116_0_x_locator0 ^ alpha116_1_x_locator1 ^ alpha116_2_x_locator2 ^ alpha116_3_x_locator3)), (~| (alpha115_0_x_locator0 ^ alpha115_1_x_locator1 ^ alpha115_2_x_locator2 ^ alpha115_3_x_locator3)), (~| (alpha114_0_x_locator0 ^ alpha114_1_x_locator1 ^ alpha114_2_x_locator2 ^ alpha114_3_x_locator3)), (~| (alpha113_0_x_locator0 ^ alpha113_1_x_locator1 ^ alpha113_2_x_locator2 ^ alpha113_3_x_locator3)), (~| (alpha112_0_x_locator0 ^ alpha112_1_x_locator1 ^ alpha112_2_x_locator2 ^ alpha112_3_x_locator3)), (~| (alpha111_0_x_locator0 ^ alpha111_1_x_locator1 ^ alpha111_2_x_locator2 ^ alpha111_3_x_locator3)), (~| (alpha110_0_x_locator0 ^ alpha110_1_x_locator1 ^ alpha110_2_x_locator2 ^ alpha110_3_x_locator3)), (~| (alpha109_0_x_locator0 ^ alpha109_1_x_locator1 ^ alpha109_2_x_locator2 ^ alpha109_3_x_locator3)), (~| (alpha108_0_x_locator0 ^ alpha108_1_x_locator1 ^ alpha108_2_x_locator2 ^ alpha108_3_x_locator3)), (~| (alpha107_0_x_locator0 ^ alpha107_1_x_locator1 ^ alpha107_2_x_locator2 ^ alpha107_3_x_locator3)), (~| (alpha106_0_x_locator0 ^ alpha106_1_x_locator1 ^ alpha106_2_x_locator2 ^ alpha106_3_x_locator3)), (~| (alpha105_0_x_locator0 ^ alpha105_1_x_locator1 ^ alpha105_2_x_locator2 ^ alpha105_3_x_locator3)), (~| (alpha104_0_x_locator0 ^ alpha104_1_x_locator1 ^ alpha104_2_x_locator2 ^ alpha104_3_x_locator3)), (~| (alpha103_0_x_locator0 ^ alpha103_1_x_locator1 ^ alpha103_2_x_locator2 ^ alpha103_3_x_locator3)), (~| (alpha102_0_x_locator0 ^ alpha102_1_x_locator1 ^ alpha102_2_x_locator2 ^ alpha102_3_x_locator3)), (~| (alpha101_0_x_locator0 ^ alpha101_1_x_locator1 ^ alpha101_2_x_locator2 ^ alpha101_3_x_locator3)), (~| (alpha100_0_x_locator0 ^ alpha100_1_x_locator1 ^ alpha100_2_x_locator2 ^ alpha100_3_x_locator3)), (~| (alpha99_0_x_locator0 ^ alpha99_1_x_locator1 ^ alpha99_2_x_locator2 ^ alpha99_3_x_locator3)), (~| (alpha98_0_x_locator0 ^ alpha98_1_x_locator1 ^ alpha98_2_x_locator2 ^ alpha98_3_x_locator3)), (~| (alpha97_0_x_locator0 ^ alpha97_1_x_locator1 ^ alpha97_2_x_locator2 ^ alpha97_3_x_locator3)), (~| (alpha96_0_x_locator0 ^ alpha96_1_x_locator1 ^ alpha96_2_x_locator2 ^ alpha96_3_x_locator3)), (~| (alpha95_0_x_locator0 ^ alpha95_1_x_locator1 ^ alpha95_2_x_locator2 ^ alpha95_3_x_locator3)), (~| (alpha94_0_x_locator0 ^ alpha94_1_x_locator1 ^ alpha94_2_x_locator2 ^ alpha94_3_x_locator3)), (~| (alpha93_0_x_locator0 ^ alpha93_1_x_locator1 ^ alpha93_2_x_locator2 ^ alpha93_3_x_locator3)), (~| (alpha92_0_x_locator0 ^ alpha92_1_x_locator1 ^ alpha92_2_x_locator2 ^ alpha92_3_x_locator3)), (~| (alpha91_0_x_locator0 ^ alpha91_1_x_locator1 ^ alpha91_2_x_locator2 ^ alpha91_3_x_locator3)), (~| (alpha90_0_x_locator0 ^ alpha90_1_x_locator1 ^ alpha90_2_x_locator2 ^ alpha90_3_x_locator3)), (~| (alpha89_0_x_locator0 ^ alpha89_1_x_locator1 ^ alpha89_2_x_locator2 ^ alpha89_3_x_locator3)), (~| (alpha88_0_x_locator0 ^ alpha88_1_x_locator1 ^ alpha88_2_x_locator2 ^ alpha88_3_x_locator3)), (~| (alpha87_0_x_locator0 ^ alpha87_1_x_locator1 ^ alpha87_2_x_locator2 ^ alpha87_3_x_locator3)), (~| (alpha86_0_x_locator0 ^ alpha86_1_x_locator1 ^ alpha86_2_x_locator2 ^ alpha86_3_x_locator3)), (~| (alpha85_0_x_locator0 ^ alpha85_1_x_locator1 ^ alpha85_2_x_locator2 ^ alpha85_3_x_locator3)), (~| (alpha84_0_x_locator0 ^ alpha84_1_x_locator1 ^ alpha84_2_x_locator2 ^ alpha84_3_x_locator3)), (~| (alpha83_0_x_locator0 ^ alpha83_1_x_locator1 ^ alpha83_2_x_locator2 ^ alpha83_3_x_locator3)), (~| (alpha82_0_x_locator0 ^ alpha82_1_x_locator1 ^ alpha82_2_x_locator2 ^ alpha82_3_x_locator3)), (~| (alpha81_0_x_locator0 ^ alpha81_1_x_locator1 ^ alpha81_2_x_locator2 ^ alpha81_3_x_locator3)), (~| (alpha80_0_x_locator0 ^ alpha80_1_x_locator1 ^ alpha80_2_x_locator2 ^ alpha80_3_x_locator3)), (~| (alpha79_0_x_locator0 ^ alpha79_1_x_locator1 ^ alpha79_2_x_locator2 ^ alpha79_3_x_locator3)), (~| (alpha78_0_x_locator0 ^ alpha78_1_x_locator1 ^ alpha78_2_x_locator2 ^ alpha78_3_x_locator3)), (~| (alpha77_0_x_locator0 ^ alpha77_1_x_locator1 ^ alpha77_2_x_locator2 ^ alpha77_3_x_locator3)), (~| (alpha76_0_x_locator0 ^ alpha76_1_x_locator1 ^ alpha76_2_x_locator2 ^ alpha76_3_x_locator3)), (~| (alpha75_0_x_locator0 ^ alpha75_1_x_locator1 ^ alpha75_2_x_locator2 ^ alpha75_3_x_locator3)), (~| (alpha74_0_x_locator0 ^ alpha74_1_x_locator1 ^ alpha74_2_x_locator2 ^ alpha74_3_x_locator3)), (~| (alpha73_0_x_locator0 ^ alpha73_1_x_locator1 ^ alpha73_2_x_locator2 ^ alpha73_3_x_locator3)), (~| (alpha72_0_x_locator0 ^ alpha72_1_x_locator1 ^ alpha72_2_x_locator2 ^ alpha72_3_x_locator3)), (~| (alpha71_0_x_locator0 ^ alpha71_1_x_locator1 ^ alpha71_2_x_locator2 ^ alpha71_3_x_locator3)), (~| (alpha70_0_x_locator0 ^ alpha70_1_x_locator1 ^ alpha70_2_x_locator2 ^ alpha70_3_x_locator3)), (~| (alpha69_0_x_locator0 ^ alpha69_1_x_locator1 ^ alpha69_2_x_locator2 ^ alpha69_3_x_locator3)), (~| (alpha68_0_x_locator0 ^ alpha68_1_x_locator1 ^ alpha68_2_x_locator2 ^ alpha68_3_x_locator3)), (~| (alpha67_0_x_locator0 ^ alpha67_1_x_locator1 ^ alpha67_2_x_locator2 ^ alpha67_3_x_locator3)), (~| (alpha66_0_x_locator0 ^ alpha66_1_x_locator1 ^ alpha66_2_x_locator2 ^ alpha66_3_x_locator3)), (~| (alpha65_0_x_locator0 ^ alpha65_1_x_locator1 ^ alpha65_2_x_locator2 ^ alpha65_3_x_locator3)), (~| (alpha64_0_x_locator0 ^ alpha64_1_x_locator1 ^ alpha64_2_x_locator2 ^ alpha64_3_x_locator3)), (~| (alpha63_0_x_locator0 ^ alpha63_1_x_locator1 ^ alpha63_2_x_locator2 ^ alpha63_3_x_locator3)), (~| (alpha62_0_x_locator0 ^ alpha62_1_x_locator1 ^ alpha62_2_x_locator2 ^ alpha62_3_x_locator3)), (~| (alpha61_0_x_locator0 ^ alpha61_1_x_locator1 ^ alpha61_2_x_locator2 ^ alpha61_3_x_locator3)), (~| (alpha60_0_x_locator0 ^ alpha60_1_x_locator1 ^ alpha60_2_x_locator2 ^ alpha60_3_x_locator3)), (~| (alpha59_0_x_locator0 ^ alpha59_1_x_locator1 ^ alpha59_2_x_locator2 ^ alpha59_3_x_locator3)), (~| (alpha58_0_x_locator0 ^ alpha58_1_x_locator1 ^ alpha58_2_x_locator2 ^ alpha58_3_x_locator3)), (~| (alpha57_0_x_locator0 ^ alpha57_1_x_locator1 ^ alpha57_2_x_locator2 ^ alpha57_3_x_locator3)), (~| (alpha56_0_x_locator0 ^ alpha56_1_x_locator1 ^ alpha56_2_x_locator2 ^ alpha56_3_x_locator3)), (~| (alpha55_0_x_locator0 ^ alpha55_1_x_locator1 ^ alpha55_2_x_locator2 ^ alpha55_3_x_locator3)), (~| (alpha54_0_x_locator0 ^ alpha54_1_x_locator1 ^ alpha54_2_x_locator2 ^ alpha54_3_x_locator3)), (~| (alpha53_0_x_locator0 ^ alpha53_1_x_locator1 ^ alpha53_2_x_locator2 ^ alpha53_3_x_locator3)), (~| (alpha52_0_x_locator0 ^ alpha52_1_x_locator1 ^ alpha52_2_x_locator2 ^ alpha52_3_x_locator3)), (~| (alpha51_0_x_locator0 ^ alpha51_1_x_locator1 ^ alpha51_2_x_locator2 ^ alpha51_3_x_locator3)), (~| (alpha50_0_x_locator0 ^ alpha50_1_x_locator1 ^ alpha50_2_x_locator2 ^ alpha50_3_x_locator3)), (~| (alpha49_0_x_locator0 ^ alpha49_1_x_locator1 ^ alpha49_2_x_locator2 ^ alpha49_3_x_locator3)), (~| (alpha48_0_x_locator0 ^ alpha48_1_x_locator1 ^ alpha48_2_x_locator2 ^ alpha48_3_x_locator3)), (~| (alpha47_0_x_locator0 ^ alpha47_1_x_locator1 ^ alpha47_2_x_locator2 ^ alpha47_3_x_locator3)), (~| (alpha46_0_x_locator0 ^ alpha46_1_x_locator1 ^ alpha46_2_x_locator2 ^ alpha46_3_x_locator3)), (~| (alpha45_0_x_locator0 ^ alpha45_1_x_locator1 ^ alpha45_2_x_locator2 ^ alpha45_3_x_locator3)), (~| (alpha44_0_x_locator0 ^ alpha44_1_x_locator1 ^ alpha44_2_x_locator2 ^ alpha44_3_x_locator3)), (~| (alpha43_0_x_locator0 ^ alpha43_1_x_locator1 ^ alpha43_2_x_locator2 ^ alpha43_3_x_locator3)), (~| (alpha42_0_x_locator0 ^ alpha42_1_x_locator1 ^ alpha42_2_x_locator2 ^ alpha42_3_x_locator3)), (~| (alpha41_0_x_locator0 ^ alpha41_1_x_locator1 ^ alpha41_2_x_locator2 ^ alpha41_3_x_locator3)), (~| (alpha40_0_x_locator0 ^ alpha40_1_x_locator1 ^ alpha40_2_x_locator2 ^ alpha40_3_x_locator3)), (~| (alpha39_0_x_locator0 ^ alpha39_1_x_locator1 ^ alpha39_2_x_locator2 ^ alpha39_3_x_locator3)), (~| (alpha38_0_x_locator0 ^ alpha38_1_x_locator1 ^ alpha38_2_x_locator2 ^ alpha38_3_x_locator3)), (~| (alpha37_0_x_locator0 ^ alpha37_1_x_locator1 ^ alpha37_2_x_locator2 ^ alpha37_3_x_locator3)), (~| (alpha36_0_x_locator0 ^ alpha36_1_x_locator1 ^ alpha36_2_x_locator2 ^ alpha36_3_x_locator3)), (~| (alpha35_0_x_locator0 ^ alpha35_1_x_locator1 ^ alpha35_2_x_locator2 ^ alpha35_3_x_locator3)), (~| (alpha34_0_x_locator0 ^ alpha34_1_x_locator1 ^ alpha34_2_x_locator2 ^ alpha34_3_x_locator3)), (~| (alpha33_0_x_locator0 ^ alpha33_1_x_locator1 ^ alpha33_2_x_locator2 ^ alpha33_3_x_locator3)), (~| (alpha32_0_x_locator0 ^ alpha32_1_x_locator1 ^ alpha32_2_x_locator2 ^ alpha32_3_x_locator3)), (~| (alpha31_0_x_locator0 ^ alpha31_1_x_locator1 ^ alpha31_2_x_locator2 ^ alpha31_3_x_locator3)), (~| (alpha30_0_x_locator0 ^ alpha30_1_x_locator1 ^ alpha30_2_x_locator2 ^ alpha30_3_x_locator3)), (~| (alpha29_0_x_locator0 ^ alpha29_1_x_locator1 ^ alpha29_2_x_locator2 ^ alpha29_3_x_locator3)), (~| (alpha28_0_x_locator0 ^ alpha28_1_x_locator1 ^ alpha28_2_x_locator2 ^ alpha28_3_x_locator3)), (~| (alpha27_0_x_locator0 ^ alpha27_1_x_locator1 ^ alpha27_2_x_locator2 ^ alpha27_3_x_locator3)), (~| (alpha26_0_x_locator0 ^ alpha26_1_x_locator1 ^ alpha26_2_x_locator2 ^ alpha26_3_x_locator3)), (~| (alpha25_0_x_locator0 ^ alpha25_1_x_locator1 ^ alpha25_2_x_locator2 ^ alpha25_3_x_locator3)), (~| (alpha24_0_x_locator0 ^ alpha24_1_x_locator1 ^ alpha24_2_x_locator2 ^ alpha24_3_x_locator3)), (~| (alpha23_0_x_locator0 ^ alpha23_1_x_locator1 ^ alpha23_2_x_locator2 ^ alpha23_3_x_locator3)), (~| (alpha22_0_x_locator0 ^ alpha22_1_x_locator1 ^ alpha22_2_x_locator2 ^ alpha22_3_x_locator3)), (~| (alpha21_0_x_locator0 ^ alpha21_1_x_locator1 ^ alpha21_2_x_locator2 ^ alpha21_3_x_locator3)), (~| (alpha20_0_x_locator0 ^ alpha20_1_x_locator1 ^ alpha20_2_x_locator2 ^ alpha20_3_x_locator3)), (~| (alpha19_0_x_locator0 ^ alpha19_1_x_locator1 ^ alpha19_2_x_locator2 ^ alpha19_3_x_locator3)), (~| (alpha18_0_x_locator0 ^ alpha18_1_x_locator1 ^ alpha18_2_x_locator2 ^ alpha18_3_x_locator3)), (~| (alpha17_0_x_locator0 ^ alpha17_1_x_locator1 ^ alpha17_2_x_locator2 ^ alpha17_3_x_locator3)), (~| (alpha16_0_x_locator0 ^ alpha16_1_x_locator1 ^ alpha16_2_x_locator2 ^ alpha16_3_x_locator3)), (~| (alpha15_0_x_locator0 ^ alpha15_1_x_locator1 ^ alpha15_2_x_locator2 ^ alpha15_3_x_locator3)), (~| (alpha14_0_x_locator0 ^ alpha14_1_x_locator1 ^ alpha14_2_x_locator2 ^ alpha14_3_x_locator3)), (~| (alpha13_0_x_locator0 ^ alpha13_1_x_locator1 ^ alpha13_2_x_locator2 ^ alpha13_3_x_locator3)), (~| (alpha12_0_x_locator0 ^ alpha12_1_x_locator1 ^ alpha12_2_x_locator2 ^ alpha12_3_x_locator3)), (~| (alpha11_0_x_locator0 ^ alpha11_1_x_locator1 ^ alpha11_2_x_locator2 ^ alpha11_3_x_locator3)), (~| (alpha10_0_x_locator0 ^ alpha10_1_x_locator1 ^ alpha10_2_x_locator2 ^ alpha10_3_x_locator3)), (~| (alpha9_0_x_locator0 ^ alpha9_1_x_locator1 ^ alpha9_2_x_locator2 ^ alpha9_3_x_locator3)), (~| (alpha8_0_x_locator0 ^ alpha8_1_x_locator1 ^ alpha8_2_x_locator2 ^ alpha8_3_x_locator3)), (~| (alpha7_0_x_locator0 ^ alpha7_1_x_locator1 ^ alpha7_2_x_locator2 ^ alpha7_3_x_locator3)), (~| (alpha6_0_x_locator0 ^ alpha6_1_x_locator1 ^ alpha6_2_x_locator2 ^ alpha6_3_x_locator3)), (~| (alpha5_0_x_locator0 ^ alpha5_1_x_locator1 ^ alpha5_2_x_locator2 ^ alpha5_3_x_locator3)), (~| (alpha4_0_x_locator0 ^ alpha4_1_x_locator1 ^ alpha4_2_x_locator2 ^ alpha4_3_x_locator3)), (~| (alpha3_0_x_locator0 ^ alpha3_1_x_locator1 ^ alpha3_2_x_locator2 ^ alpha3_3_x_locator3)), (~| (alpha2_0_x_locator0 ^ alpha2_1_x_locator1 ^ alpha2_2_x_locator2 ^ alpha2_3_x_locator3)), (~| (alpha1_0_x_locator0 ^ alpha1_1_x_locator1 ^ alpha1_2_x_locator2 ^ alpha1_3_x_locator3)), (~| (alpha0_0_x_locator0 ^ alpha0_1_x_locator1 ^ alpha0_2_x_locator2 ^ alpha0_3_x_locator3))};;
endmodule

