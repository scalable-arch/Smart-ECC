module bch_ibm(syndrome1, syndrome2, syndrome3, locator0, locator1, locator2);
  input [3:0] syndrome1;
  input [3:0] syndrome2;
  input [3:0] syndrome3;
  output [3:0] locator0;
  output [3:0] locator1;
  output [3:0] locator2;

  wire [3:0] nu0_0;
  wire [3:0] nu0_1;
  wire [3:0] nu0_2;
  wire [3:0] nu2_0;
  wire [3:0] nu2_1;
  wire [3:0] nu2_2;
  wire [3:0] nu4_0;
  wire [3:0] nu4_1;
  wire [3:0] nu4_2;
  wire [3:0] kappa0_0;
  wire [3:0] kappa0_1;
  wire [3:0] kappa0_2;
  wire [3:0] kappa2_0;
  wire [3:0] kappa2_1;
  wire [3:0] kappa2_2;
  wire [3:0] kappa4_0;
  wire [3:0] kappa4_1;
  wire [3:0] kappa4_2;
  wire [3:0] delta0;
  wire [3:0] delta2;
  wire [3:0] d0;
  wire [3:0] d2;
  wire [3:0] delta0_x_nu2_0;
  wire [3:0] delta0_x_nu2_1;
  wire [3:0] delta0_x_nu2_2;
  wire [3:0] d0_x_kappa0_0;
  wire [3:0] d0_x_kappa0_1;
  wire [3:0] d0_x_kappa0_2;
  wire [3:0] d2_x_kappa2_0;
  wire [3:0] d2_x_kappa2_1;
  wire [3:0] d2_x_kappa2_2;
  wire [3:0] nu0_0_x_syndrome1;
  wire [3:0] nu2_0_x_syndrome3;
  wire [3:0] nu2_1_x_syndrome2;
  wire [3:0] nu2_2_x_syndrome1;
  wire cond0;
  wire cond2;

  gfmult gfm_delta0_x_nu2_0(delta0, nu2_0, delta0_x_nu2_0);
  gfmult gfm_delta0_x_nu2_1(delta0, nu2_1, delta0_x_nu2_1);
  gfmult gfm_delta0_x_nu2_2(delta0, nu2_2, delta0_x_nu2_2);
  gfmult gfm_d0_x_kappa0_0(d0, kappa0_0, d0_x_kappa0_0);
  gfmult gfm_d0_x_kappa0_1(d0, kappa0_1, d0_x_kappa0_1);
  gfmult gfm_d0_x_kappa0_2(d0, kappa0_2, d0_x_kappa0_2);
  gfmult gfm_d2_x_kappa2_0(d2, kappa2_0, d2_x_kappa2_0);
  gfmult gfm_d2_x_kappa2_1(d2, kappa2_1, d2_x_kappa2_1);
  gfmult gfm_d2_x_kappa2_2(d2, kappa2_2, d2_x_kappa2_2);
  gfmult gfm_nu0_0_x_syndrome1(nu0_0, syndrome1, nu0_0_x_syndrome1);
  gfmult gfm_nu2_0_x_syndrome3(nu2_0, syndrome3, nu2_0_x_syndrome3);
  gfmult gfm_nu2_1_x_syndrome2(nu2_1, syndrome2, nu2_1_x_syndrome2);
  gfmult gfm_nu2_2_x_syndrome1(nu2_2, syndrome1, nu2_2_x_syndrome1);

  assign locator0 = nu4_0;
  assign locator1 = nu4_1;
  assign locator2 = nu4_2;
  assign nu0_0 = 4'b0001;
  assign nu0_1 = 4'b0;
  assign nu0_2 = 4'b0;
  assign nu2_0 = nu0_0;
  assign nu2_1 = nu0_1 ^ d0_x_kappa0_0;
  assign nu2_2 = nu0_2 ^ d0_x_kappa0_1;
  assign nu4_0 = delta0_x_nu2_0;
  assign nu4_1 = delta0_x_nu2_1 ^ d2_x_kappa2_0;
  assign nu4_2 = delta0_x_nu2_2 ^ d2_x_kappa2_1;
  assign kappa0_0 = 4'b0001;
  assign kappa0_1 = 4'b0;
  assign kappa0_2 = 4'b0;
  assign kappa2_0 = cond0 ? 4'b0 : 4'b0;
  assign kappa2_1 = cond0 ? 4'b0 : nu0_0;
  assign kappa2_2 = cond0 ? kappa0_0 : nu0_1;
  assign kappa4_0 = cond2 ? 4'b0 : 4'b0;
  assign kappa4_1 = cond2 ? 4'b0 : nu2_0;
  assign kappa4_2 = cond2 ? kappa2_0 : nu2_1;
  assign delta0 = cond0 ? 4'b0001 : d0;
  assign delta2 = cond2 ? delta0 : d2;
  assign d0 = nu0_0_x_syndrome1 ^ nu0_1;
  assign d2 = nu2_0_x_syndrome3 ^ nu2_1_x_syndrome2 ^ nu2_2_x_syndrome1;
  assign cond0 = (~| d0) | (| nu0_1) | (| nu0_2);
  assign cond2 = (~| d2) | (| nu2_2);
endmodule
