module gfmult(a, b, c);
  input [9:0] a;
  input [9:0] b;
  output [9:0] c;

  assign c = ({10{b[0]}} & ((a << 0))) ^ ({10{b[1]}} & ((a << 1) ^ ({10{a[9]}} & 10'b0000001001))) ^ ({10{b[2]}} & ((a << 2) ^ ({10{a[9]}} & 10'b0000010010) ^ ({10{a[8]}} & 10'b0000001001))) ^ ({10{b[3]}} & ((a << 3) ^ ({10{a[9]}} & 10'b0000100100) ^ ({10{a[8]}} & 10'b0000010010) ^ ({10{a[7]}} & 10'b0000001001))) ^ ({10{b[4]}} & ((a << 4) ^ ({10{a[9]}} & 10'b0001001000) ^ ({10{a[8]}} & 10'b0000100100) ^ ({10{a[7]}} & 10'b0000010010) ^ ({10{a[6]}} & 10'b0000001001))) ^ ({10{b[5]}} & ((a << 5) ^ ({10{a[9]}} & 10'b0010010000) ^ ({10{a[8]}} & 10'b0001001000) ^ ({10{a[7]}} & 10'b0000100100) ^ ({10{a[6]}} & 10'b0000010010) ^ ({10{a[5]}} & 10'b0000001001))) ^ ({10{b[6]}} & ((a << 6) ^ ({10{a[9]}} & 10'b0100100000) ^ ({10{a[8]}} & 10'b0010010000) ^ ({10{a[7]}} & 10'b0001001000) ^ ({10{a[6]}} & 10'b0000100100) ^ ({10{a[5]}} & 10'b0000010010) ^ ({10{a[4]}} & 10'b0000001001))) ^ ({10{b[7]}} & ((a << 7) ^ ({10{a[9]}} & 10'b1001000000) ^ ({10{a[8]}} & 10'b0100100000) ^ ({10{a[7]}} & 10'b0010010000) ^ ({10{a[6]}} & 10'b0001001000) ^ ({10{a[5]}} & 10'b0000100100) ^ ({10{a[4]}} & 10'b0000010010) ^ ({10{a[3]}} & 10'b0000001001))) ^ ({10{b[8]}} & ((a << 8) ^ ({10{a[9]}} & 10'b0010001001) ^ ({10{a[8]}} & 10'b1001000000) ^ ({10{a[7]}} & 10'b0100100000) ^ ({10{a[6]}} & 10'b0010010000) ^ ({10{a[5]}} & 10'b0001001000) ^ ({10{a[4]}} & 10'b0000100100) ^ ({10{a[3]}} & 10'b0000010010) ^ ({10{a[2]}} & 10'b0000001001))) ^ ({10{b[9]}} & ((a << 9) ^ ({10{a[9]}} & 10'b0100010010) ^ ({10{a[8]}} & 10'b0010001001) ^ ({10{a[7]}} & 10'b1001000000) ^ ({10{a[6]}} & 10'b0100100000) ^ ({10{a[5]}} & 10'b0010010000) ^ ({10{a[4]}} & 10'b0001001000) ^ ({10{a[3]}} & 10'b0000100100) ^ ({10{a[2]}} & 10'b0000010010) ^ ({10{a[1]}} & 10'b0000001001)));
endmodule
