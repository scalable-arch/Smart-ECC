module SEC_encoder(input [127:0] message, output [135:0] codeword);

	assign codeword[135:8] = message[127:0];
	assign codeword[7] = ^(message&128'b01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101);
	assign codeword[6] = ^(message&128'b00110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011);
	assign codeword[5] = ^(message&128'b00001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111);
	assign codeword[4] = ^(message&128'b11111111000000001111111100000000000000001111111111111111000000001111111100000000000000001111111111111111000000000000000011111111);
	assign codeword[3] = ^(message&128'b11111111000000000000000011111111111111110000000011111111000000000000000011111111111111110000000011111111000000000000000011111111);
	assign codeword[2] = ^(message&128'b00000000111111111111111100000000111111110000000011111111000000000000000011111111000000001111111100000000111111111111111100000000);
	assign codeword[1] = ^(message&128'b00000000111111110000000011111111000000001111111100000000111111111111111100000000111111110000000011111111000000001111111100000000);
	assign codeword[0] = ^(message&128'b00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111);

endmodule
