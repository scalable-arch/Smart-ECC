module decoder_tb;
  reg [541:0] received;
  wire [541:0] codeword;
  wire [511:0] message;
  wire detection;
  integer failures;

  bch_decoder decoder(received, codeword, message, detection);

  initial
  begin
    failures = 0;

    received <= 542'b01100111000011010100011100110001001011010110100111101101001011110100110110101001001001000011001100101000011100000110000100100100011011110100011111000010000011001101010100111111111100011110010110011000001111011011010000000110011110110000010011001111000111001010001000001100011101001111111111110111101100111001110000111011111011010100011110111000110001110110001011111110111000111000011100111000001011111011100010010011001101011010101100001010001011011010111101101010111000111111100010110001101111100000101100101010000110011111010011010111000011;
    #1;
    if (message != 512'b01100111000011010100011100110001001011010110100111101101001011110100110110101001001001000011001100101000011100000110000100100100011011110100011111000010000011001101010100111111111100011110010110011000001111011011010000000110011110110000010011001111000111001010001000001100011101001111111111110111101100111001110000111011111011010100011110111000110001110110001011111110111000111000011100111000001011111011100010010011001101011010101100001010001011011010111101101010111000111111100010110001101111100000101100101010 || detection)
      failures = failures+1;

    received <= 542'b11111110111001001110110100000111110111100010000111110001001111100011110100100101010000010110000001101101000000100000101100011101000010011010001111011000010000101010001111000100001111100111101100011101000100111000101001001111111001010001111011011000001001100001010000000111110011100000111001111011000001000000101111001010100110110111000011010100111111011111101001010000000000110000000111100001110101000111101010000001100011010001011110110000111111110110100101101101011101111101011001000111010111101011011111000000100100100111000001011010111101;
    #1;
    if (message != 512'b11111110111001001110110100000111110111100010000111110001001111100011110100100101010000010110000001101101000000100000101100011101000010011010001111011000010000101010001111000100001111100111101100011101000100111000101001001111111001010001111011011000001001100001010000000111110011100000111001111011000001000000101111001010100110110111000011010100111111011111101001010000000000110000000111100001110101000111101010000001100011010001011110110000111111110110100101101101011101111101011001000111010111101011011111000000 || detection)
      failures = failures+1;

    received <= 542'b11011010111110000110011100111010001000000101011110010001110111001000000011010011010010111000100100111110111101110010101111110100111000001000101101011000011100010011111110111001111101011101101100000001011101000100011101001110100100011001110011001110010011010000110010011111100100010000011000000011011001111010110010111001101101000001110010011111111111100100110111010000111001100110100001010001001000011010110010011010001110001101000000001010110100001101111001110110001001100000011100000011110100010100000010011101101001110010101100001011001111;
    #1;
    if (message != 512'b11011010111110000110011100111010001000000101011110010001110111001000000011010011010010111000100100111110111101110010101111110100111000001000101101011000011100010011111110111001111101011101101100000001011101000100011101001110100100011001110011001110010011010000110010011111100100010000011000000011011001111010110010111001101101000001110010011111111111100100110111010000111001100110100001010001001000011010110010011010001110001101000000001010110100001101111001110110001001100000011100000011110100010100000010011101 || detection)
      failures = failures+1;

    received <= 542'b00001100011011111101000111101101000000100011010010000000010100110000011000110001111010001111000000000100001011101010000111110100110100100100100010111000010110000010011001101001001001100001110100111100010110000010100000110111100001110110100001000010000101110111111010111011110011100110111110001000001001001111001101000011100101010001111001110110010110011100001111101011100000011000000110111011111010101001110001101100010101010110011010011011011010001101100110000110010100010000011010001010101100011000011010101101101001001111110101010111100110;
    #1;
    if (message != 512'b00001100011011111101000111101101000000100011010010000000010100110000011000110001111010001111000000000100001011101010000111110100110100100100100010111000010110000010011001101001001001100001110100111100010110000010100000110111100001110110100001000010000101110111111010111011110011100110111110001000001001001111001101000011100101010001111001110110010110011100001111101011100000011000000110111011111010101001110001101100010101010110011010011011011010001101100110000110010100010000011010001010101100011000011010101101 || detection)
      failures = failures+1;

    received <= 542'b10010111001010001110101101001110101011100011101110010011011011000011001011101010000001111001110111111000000101000010001111110111101001010110000001100100110100111110101101110100100100011001000000000010100101110111110111010010101101000100101111100000101111000111100110110011111010111010110011000111101011001100111000011100100100000101010100010000001111110011101111000011001000100110100000000110111101101010011001011110000101100010101010101110011000110111011101111110111001111011110100011010101111110100110110001111100011111001100111000000110100;
    #1;
    if (message != 512'b10010111001010001110101101001110101011100011101110010011011011000011001011101010000001111001110111111000000101000010001111110111101001010110000001100100110100111110101101110100100100011001000000000010100101110111110111010010101101000100101111100000101111000111100110110011111010111010110011000111101011001100111000011100100100000101010100010000001111110011101111000011001000100110100000000110111101101010011001011110000101100010101010101110011000110111011101111110111001111011110100011010101111110100110110001111 || detection)
      failures = failures+1;

    received <= 542'b11111100010000001111011000010101101100100111110101010010000111000010011110101010100101101101011001011110111000111100101101100110110110001001110011011101010101111001100011111001110010000001001110100010011100010111110111101010101000101001001010111101000000111011001001011011000001111001010010001100111010111101001000001110101001001000000000101101011100110101100110100011001011001000011100001101111110001010000001100110000111001111100111001000010010101001001011100101001010000111110010101001101111011110110101111000101010010010111101000100111010;
    #1;
    if (message != 512'b11111100010000001111011000010101101100100111110101010010000111000010011110101010100101101101011001011110111000111100101101100110110110001001110011011101010101111001100011111001110010000001001110100010011100010111110111101010101000101001001010111101000000111011001001011011000001111001010010001100111010111101001000001110101001001000000000101101011100110101100110100011001011001000011100001101111110001010000001100110000111001111100111001000010010101001001011100101001010000111110010101001101111011110110101111000 || detection)
      failures = failures+1;

    received <= 542'b01011100011000111110001001010011100010100001101100001101010011101001011001001111111110010000111001110100001100110001101001111010111110001011100100101000010100001011101000010000100011111000111010010001000110101001000100101010011110011100001000001010000111001110000101111011010111010000010110011000111111011100111110100111001101110001110110000111010101101111110010110010000100111111110110100111001100011001110001111110000110010001011001101001111110111001110011101010100000101100011101111010010011110101010101101110110101101000100011000011001100;
    #1;
    if (message != 512'b01011100011000111110001001010011100010100001101100001101010011101001011001001111111110010000111001110100001100110001101001111010111110001011100100101000010100001011101000010000100011111000111010010001000110101001000100101010011110011100001000001010000111001110000101111011010111010000010110011000111111011100111110100111001101110001110110000111010101101111110010110010000100111111110110100111001100011001110001111110000110010001011001101001111110111001110011101010100000101100011101111010010011110101010101101110 || detection)
      failures = failures+1;

    received <= 542'b01111100111011100000000111000101010110100111011100011010000010100011000011111011011111110101101011011001011110111101111110111011101000110010101110000111111110010010110100001100011110010001000111001000001011110111101000000100101000111010101000100110100011111001110000011111010100000111000011100011101011010101000010101100001101010100111111111100000101000010100111111101001101111011100000001010001011011111101001011011110011010010001100111110011011110001011110001101110101000010010101010100110100110000101100111011101100000011000101100110011111;
    #1;
    if (message != 512'b01111100111011100000000111000101010110100111011100011010000010100011000011111011011111110101101011011001011110111101111110111011101000110010101110000111111110010010110100001100011110010001000111001000001011110111101000000100101000111010101000100110100011111001110000011111010100000111000011100011101011010101000010101100001101010100111111111100000101000010100111111101001101111011100000001010001011011111101001011011110011010010001100111110011011110001011110001101110101000010010101010100110100110000101100111011 || detection)
      failures = failures+1;

    received <= 542'b00010000000110011000101110000101011100110110110001101001000110001000011000010010011111100110000001101111110111010000100101011100000111001110000100011010011010001100010010100111110010101101011100011000101011110011111011010000101010111011100000000010010110001111000110000000001000100111001011101101101111000111111110001000010100100100001111001001000000011101111011110000000001010111011101111011101000110010100000010110100000100111101101000000110110110001100010000111101101101010110100100001100111110000100010101010110100001001001001010100101011;
    #1;
    if (message != 512'b00010000000110011000101110000101011100110110110001101001000110001000011000010010011111100110000001101111110111010000100101011100000111001110000100011010011010001100010010100111110010101101011100011000101011110011111011010000101010111011100000000010010110001111000110000000001000100111001011101101101111000111111110001000010100100100001111001001000000011101111011110000000001010111011101111011101000110010100000010110100000100111101101000000110110110001100010000111101101101010110100100001100111110000100010101010 || detection)
      failures = failures+1;

    received <= 542'b00000110111001111100110100110001111001110100110000111011100101110010011011111011010001101100000000101011010110001110000001010101100000111001000101011100011011000111110110001011111100100010010111110010001111010111010000111101101001001000110000000110001010111110000111100110010111011011011110111101010111000011100000000011010000101001010100001010010010101110011111010101111110001011011101000011010001101100101101111000001011110111100011000111101111011001000010101111000111001101010110110111110001110001011011100001100111111010010100000100010101;
    #1;
    if (message != 512'b00000110111001111100110100110001111001110100110000111011100101110010011011111011010001101100000000101011010110001110000001010101100000111001000101011100011011000111110110001011111100100010010111110010001111010111010000111101101001001000110000000110001010111110000111100110010111011011011110111101010111000011100000000011010000101001010100001010010010101110011111010101111110001011011101000011010001101100101101111000001011110111100011000111101111011001000010101111000111001101010110110111110001110001011011100001 || detection)
      failures = failures+1;

    received <= 542'b11001010001000100110111100000011110010001000110001001001000111101101000101001001000111111110100001001011001111111010000010000000000111010001011001100110000101100111110001011000010101000111001001000100110001010100111111111111100110010101101011011111100111010001101001011100011010010100011000110111100000100010101010100000011101110001100011101001101110111000000111111001100100101011111001001000111001111001111101110101010101010000111000110000110001110100001000010010100001110011011000110010111010010100111010000110110001110110110100011010110101;
    #1;
    if (message != 512'b11001010001000100110111100000011110010001000110001001001000111101101000101001001000111111110100001001011001111111010000010000000000111010001011001100110000101100111110001011000010101000111001001000100110001010100111111111111100110010101101011011111100111010001101001011100011010010100011000110111100000100010101010100000011101110001100011101001101110111000000111111001100100101011111001001000111001111001111101110101010101010000111000110000110001110100001000010010100001110011011000110010111010010100111010000110 || detection)
      failures = failures+1;

    received <= 542'b11001100110111011000111110101011101000110010111000101010101011110111010011101001010001110001110011010111010101001110101111011110111001101011100011100000101101100101111111101110010010101101100011111001011011101111100100010000100111001000101000110110000111011000111010111101000001010001111111001001000011001111110111101101111001110011110110000001100110100001001011000101001101001011011110100000111100000100001000001110101001111110011011000101011110011111110100110111101100110000000000101001101100000000101110101101100011000100101001011101101111;
    #1;
    if (message != 512'b11001100110111011000111110101011101000110010111000101010101011110111010011101001010001110001110011010111010101001110101111011110111001101011100011100000101101100101111111101110010010101101100011111001011011101111100100010000100111001000101000110110000111011000111010111101000001010001111111001001000011001111110111101101111001110011110110000001100110100001001011000101001101001011011110100000111100000100001000001110101001111110011011000101011110011111110100110111101100110000000000101001101100000000101110101101 || detection)
      failures = failures+1;

    received <= 542'b11011000111110111111101100001111100110000010011000000011110110101010000100101010001001001011001100111011110001110101110110001000100110000101110011011101010011000000000010001111010011001100111100001101110011000110010100000011010110000010100010001001110000111111110100110111010111001001110100010010000111001000110010110111100011001110011101110011001110001110101010001100111001011001101101010011010011101110010011011110010110000101100011001101011001101010010100101100011010100001001001011100010011001110111100010001100100110011111000111000100011;
    #1;
    if (message != 512'b11011000111110111111101100001111100110000010011000000011110110101010000100101010001001001011001100111011110001110101110110001000100110000101110011011101010011000000000010001111010011001100111100001101110011000110010100000011010110000010100010001001110000111111110100110111010111001001110100010010000111001000110010110111100011001110011101110011001110001110101010001100111001011001101101010011010011101110010011011110010110000101100011001101011001101010010100101100011010100001001001011100010011001110111100010001 || detection)
      failures = failures+1;

    received <= 542'b10100000000111011111101111001100000010111101100000000000001100111101000000000111100011000001101110101100010001011011110110001100101011011111001010001001011111111110001010111010100111110010111000110000110110011001010000011000011011000011011111100010100011111010011101111010001100101010100101110001011110111011111001101001010110110101011010111111101110100110101010010111001011010101011010011111001010110111000000000110010101100101001110101000101110100101000001010001001001010110000111111000011110100000000101100011100110011111010101110110101100;
    #1;
    if (message != 512'b10100000000111011111101111001100000010111101100000000000001100111101000000000111100011000001101110101100010001011011110110001100101011011111001010001001011111111110001010111010100111110010111000110000110110011001010000011000011011000011011111100010100011111010011101111010001100101010100101110001011110111011111001101001010110110101011010111111101110100110101010010111001011010101011010011111001010110111000000000110010101100101001110101000101110100101000001010001001001010110000111111000011110100000000101100011 || detection)
      failures = failures+1;

    received <= 542'b00000101010100011100011110000101010100001010101000111010101111100100010000101011000010100110010101111100000111000101000000011111001100001110011111110101011101111001101100100110101100001011000000000111100011101101000101111110111110111010110010011010011010111100010110111001111000111100011101010101101001011100110000101111000010111101011010101100011101101000001111011001011011101011110011010000110101011101010101011101011100010010110100011101001001101111010010000011101010010000011100011001101110010000001001001111000010100000110100011001110110;
    #1;
    if (message != 512'b00000101010100011100011110000101010100001010101000111010101111100100010000101011000010100110010101111100000111000101000000011111001100001110011111110101011101111001101100100110101100001011000000000111100011101101000101111110111110111010110010011010011010111100010110111001111000111100011101010101101001011100110000101111000010111101011010101100011101101000001111011001011011101011110011010000110101011101010101011101011100010010110100011101001001101111010010000011101010010000011100011001101110010000001001001111 || detection)
      failures = failures+1;

    received <= 542'b10100111001100010100101100111001110000001010100001100110101001110010100001000010100011111111001101101100111011101110001001100001101010111100110011000001110111010101010010101101111111001000001111011100001101101111010110111111111101010000001100111001011000010001110100011011100001011110111101000001111101010110000101000000111011001011010110100010101100000111001111011110000111110111101011101000001101100100011000010001100110001101001000100100101011001101111011101100001011100111010100110011010101100100101010011000010011111111111111111111011101;
    #1;
    if (message != 512'b10100111001100010100101100111001110000001010100001100110101001110010100001000010100011111111001101101100111011101110001001100001101010111100110011000001110111010101010010101101111111001000001111011100001101101111010110111111111101010000001100111001011000010001110100011011100001011110111101000001111101010110000101000000111011001011010110100010101100000111001111011110000111110111101011101000001101100100011000010001100110001101001000100100101011001101111011101100001011100111010100110011010101100100101010011000 || detection)
      failures = failures+1;

    received <= 542'b10101110111111000001011001101111100111010001001011110110111100000100011000011111110010101100010100011101001000010100110110000101000110100110101111110110111110110001011000101010100111101111100101011000011100100110010000111100010010011100110000011110110101101111001110011101110011000100000011110000000001010000010001001110111000011110011010001111110110010101000011100101011110001111010101111100011110101010110100110111000000111010011011001111111000000010001010101011111010010001101000010111001110101100110100001100011110111010101001110100011011;
    #1;
    if (message != 512'b10101110111111000001011001101111100111010001001011110110111100000100011000011111110010101100010100011101001000010100110110000101000110100110101111110110111110110001011000101010100111101111100101011000011100100110010000111100010010011100110000011110110101101111001110011101110011000100000011110000000001010000010001001110111000011110011010001111110110010101000011100101011110001111010101111100011110101010110100110111000000111010011011001111111000000010001010101011111010010001101000010111001110101100110100001100 || detection)
      failures = failures+1;

    received <= 542'b10000100001000111100011100011110011000001001101110001110101010001100010101011111111001011101100111011010010011111110000010101101111000010010011111001011111000010001101111101010011110111110010001110111110100011110100001101010000100001110101111001111010010000110011011001100011100011011011011001100111011110000111111001001010011010111110010000100010101101000111011100001101100011001101111001101101000011000010010010100010110010111101000100000101010000101111001000010101010110110110010011001101000010011111111001100111011100001000000010010100001;
    #1;
    if (message != 512'b10000100001000111100011100011110011000001001101110001110101010001100010101011111111001011101100111011010010011111110000010101101111000010010011111001011111000010001101111101010011110111110010001110111110100011110100001101010000100001110101111001111010010000110011011001100011100011011011011001100111011110000111111001001010011010111110010000100010101101000111011100001101100011001101111001101101000011000010010010100010110010111101000100000101010000101111001000010101010110110110010011001101000010011111111001100 || detection)
      failures = failures+1;

    received <= 542'b01101111100001101111110011111100000101110011000011010010000001010010111101101011110001101100011011000110110101100001110010100100111100110001111010011110011101010001101001000010000000101110100110100100111010101010000000000100010111101011010010001010000001100110010110110101001101111011000110100111000110010100000000000110001011110110001001011100010101000111011101001110010000000111010101101001010111010101001111010111101110010101101110011001011011011101001001100110010000101101011010011011101111111111000101001111110001000001101110100011001001;
    #1;
    if (message != 512'b01101111100001101111110011111100000101110011000011010010000001010010111101101011110001101100011011000110110101100001110010100100111100110001111010011110011101010001101001000010000000101110100110100100111010101010000000000100010111101011010010001010000001100110010110110101001101111011000110100111000110010100000000000110001011110110001001011100010101000111011101001110010000000111010101101001010111010101001111010111101110010101101110011001011011011101001001100110010000101101011010011011101111111111000101001111 || detection)
      failures = failures+1;

    received <= 542'b01000110011001111001111101101001000011001100011000010001100100001001010010110001110010101010100101001100001110010111010101010000101001100011111111111001001010100001101001101100001100111110010010110100001110011101101110000111110011010011000100010001000100101011101101000001100010011011101001110101000011111000101111000011100010100100111011011111010011011010110001001101000001100100001010010001101000000111001001010001000101000000100010110010110110010010101101010111010101011000000001111110000100111111001111101010101111110101011000000010000011;
    #1;
    if (message != 512'b01000110011001111001111101101001000011001100011000010001100100001001010010110001110010101010100101001100001110010111010101010000101001100011111111111001001010100001101001101100001100111110010010110100001110011101101110000111110011010011000100010001000100101011101101000001100010011011101001110101000011111000101111000011100010100100111011011111010011011010110001001101000001100100001010010001101000000111001001010001000101000000100010110010110110010010101101010111010101011000000001111110000100111111001111101010 || detection)
      failures = failures+1;

    received <= 542'b11001000111010001110101100100000101101001100100100010010100111110011011100000101011001111110100110000000001101101000111010100110111110000110110010111011000110101101001110110000100101000110101001111000001000000101001001110101010010000110110011101100001110101000011000011100110011001101110010000010001000111110101001010010100011110010111010011101101000110000010100011111001110000000111110000100111101010110001110000111110101011110001000101001000111110001010100111101000001110011011001010000000101001000011010000101010110101110101000111010011010;
    #1;
    if (message != 512'b11001000111010001110101100100000101101001100100100010010100111110011011100000101011001111110100110000000001101101000111010100110111110000110110010111011000110101101001110110000100101000110101001111000001000000101001001110101010010000110110011101100001110101000011000011100110011001101110010000010001000111110101001010010100011110010111010001101101000110000010100011111001110000000111110000100111101010110001110000111110101011110001000101001000111110001010100111101000001110011011001010000000101001000011010000101 || !detection)
      failures = failures+1;

    received <= 542'b11001100100001111010001001111010110111001110110010001101111010001010110101010111010101001100010000101101110111100000010001110000001001011101011100111111000001101101100101111000010100011011110110110010010010000100101111001001000100011101010001001010011000111101110011110000010111111001100001101001100110011001001011010011111101011100010010110101001011000010100010100101110010011101011111101001000111000111111011011001011100010001100000001111000000011110111101110000010010111110110000100000111001110110000000101000001011001110000001011101101100;
    #1;
    if (message != 512'b11001100100001111010001001111010110111001110110010001101111010001010110101010111010101001100010000101101110111100000010001110000001001011101011100111111000001101101100101111000010100011011110110110010010010000100101110001001000100011101010001001010011000111101110011110000010111111001100001101001100110011001001011010011111101011100010010110101001011000010100010100101110010011101011111101001000111000111111011011001011100010001100000001111000000011110111101110000010010111110110000100000111001110110000000101000 || !detection)
      failures = failures+1;

    received <= 542'b11101001101110100111100101101010100111011100011111010101000111110100110111111001011000011010000100000111100010000010001101111101100001010101101111111011001101010110001111000100101101111111110101100011001110010110100100111011110111000100111111000011000000000000001100111010110011010100010101100001000011010010110001111101110110101101110010011010100011101010001011111000100100110101001111111011001111100000110100010100101111110000111111100101101100011100000110101011011101100001100111001101100001001010101010101010111101100100010110100110100001;
    #1;
    if (message != 512'b11101001101110100111100101101010100111011100011111010101000111110100110111111001011000011010000100000111100010000010001101111101100001010101101111111011001101010110001111000100101101111111110101100011001110010110100100111011110111000100111111000011000000000000001100111010110011010100010101100001000011010010110001111101110110100101110010011010100011101010001011111000100100110101001111111011001111100000110100010100101111110000111111100101101100011100000110101011011101100001100111001101100001001010101010101010 || !detection)
      failures = failures+1;

    received <= 542'b01101000100000011101011010100110000101101000001111010000011111001000011000101100110011010010110011101000000011011001111001101101100010010011100001100100011001011010111101000111101101110100010110100101011101110100101000100010000101111111110011000010001001100001111000110010010101010101011101110100111001101000000011100111101110010100010110010110011110001100001000101111101100100100000011110001111000110100110000011011011111110010110101010010010010001100001100111101000011101110011011001110010001100100000110100001111000010010101000000011100111;
    #1;
    if (message != 512'b01101000100000011101011010100110000101101000001111010000011111001000011000101100110011010010110011101000000011011001111001101101100010010011100001100100011001011010111101000111101101110100010110100101011101110100101000100010000101111111110011000010001001100001111000110010010101010101011101110100111001001000000011100111101110010100010110010110011110001100001000101111101100100100000011110001111000110100110000011011011111110010110101010010010010001100001100111101000011101110011011001110010001100100000110100001 || !detection)
      failures = failures+1;

    received <= 542'b11011100100001010011011001100111110010111111100001010001000000011101000011111111110000001110100101110111110001011001101011001010001001001101011000111110000001100001001101101110000000110111100000101011100010011010110001000001000101001111000011110110110010000000001011100101001011101011100001111010111111000010111100000110011101100100000001001110010011101100101010001001001001101010000100100110000100111000011111111011111111010110111001001000111111110001010010010001100100100110001110100000111101100000001100010011000100100000011111110101001110;
    #1;
    if (message != 512'b11011100100001000011011001100111110010111111100001010001000000011101000011111111110000001110100101110111110001011001101011001010001001001101011000111110000001100001001101101110000000110111100000101011100010011010110001000001000101001111000011110110110010000000001011100101001011101011100001111010111111000010111100000110011101100100000001001110010011101100101010001001001001101010000100100110000100111000011111111011111111010110111001001000111111110001010010010001100100100110001110100000111101100000001100010011 || !detection)
      failures = failures+1;

    received <= 542'b01101001100011010001011000010011110011111100100111101011001000011010101101111110101001000111000000010011100010001101101011111010001001010001100111111000001000110101010110000111011010010000010110011110100010110111001010010100100000101101010111001100110000010100011001100100111011011011111110101011111000101111000111001100110100011001101011111011111010101011011101011101100010110101111111110011000011001110010001111100011010001001001100010101111110001001000100000011000010100111011000001001011111001111010011111010111000011110110101010100011010;
    #1;
    if (message != 512'b01101001100011010001011000010011110011111100100111101011001000011010101101111110101001000111000000010011100010001101101011111010001001010001100111111000001000110101010110001111011010010000010110011110100010110111001010010100100000101101010111001100110000010100011001100100111011011011111110101011111000101111000111001100110100011001101011111011111010101011011101011101100010110101111111110011000011001110010001111100011010001001001100010101111110001001000100000011000010100111011000001001011111001111010011111010 || !detection)
      failures = failures+1;

    received <= 542'b10011011111101101001000010001110000110011111110011010101110000101110100011101010001110111001001110010111101001110001101110010000010011100110110110100110001111001000110111011101110110010101110110001000010100010001101000000001000011100010110100001000000001011000011100000001110100110011111000001000110001001100000001100110010101111110001100101110000010011100011001000100011000110001000100111101000011101011000111110001001110111111001101010100101101101100010101011100111111001110010000001001111001010011100011101001000000011000011100000111111000;
    #1;
    if (message != 512'b10011011111101101001000010001110000110011111110011010101110000101110100011101010001110111001001110010111101001110001101110010000010011100110110110100110001111001000110111011101110110010101110110001000010100010001101000000001000011100010110100001000000001011000011100000001110100110011111000001000110001001100000001100110010101111110001100101110000010011100011001000100011000110001000100111101000011101011000111110001001110111111001101010100101101101100010101011100111111001110010000011001111001010011100011101001 || !detection)
      failures = failures+1;

    received <= 542'b01011111110001111010110110000101000111010110111111000111101110001010101000010100010100111111101011101011110111011111011101100010010001010000110011001000101111101100001000101100011100011101111101100100100101101111101111101010000000100110101110001101101100110000101000110011000101111111101110101010100001100111001011100110000001000111001011011010101100111110001110011000111001000001000010001001010110100110100111001000000010001111110001111100011100101000100010010101111010011111101001000000000010110011010110100111100111110011101110101011000111;
    #1;
    if (message != 512'b01011111110001111010110110000101000111010110111111000111101110001010101000010100010100111111101011101011110111011111011101100010010001010000110011001000101111101100001000101100011100011101111101100100100101101111101111101010000000100110101110001101101100110000101000110011000101111111101110101010100001100111001011100110000001000111001011011010101100111110001110011000111001000001000010001001010110100110100111001000000010001111110001111100011100101100100010010101111010011111101001000000000010110011010110100111 || !detection)
      failures = failures+1;

    received <= 542'b00100101010100010001011110101111000111001101001000110101111010110110110001101111011001001010100100010001100010000101100111110111111010100000010001100100010111110010100110100001001111011101010010000100011100100010101101001001010011010110010100110011110000000001110111101001111001010101101001101110010111010010010110110101001001110000000000000000100000111010101001101011110001001110001010001100101101010011010000101101111011100010000001011110001111110010010001100100110100011101001000001101110010100110001001010101001101000100100010100101101010;
    #1;
    if (message != 512'b00100101010100010001011110101111000111001101001000110101111010110110110001101111011001001010100100010001100010000101100111110111111010100000010001100100010111110010100110100000001111011101010010000100011100100010101101001001010011010110010100110011110000000001110111101001111001010101101001101110010111010010010110110101001001110000000000000000100000111010101001101011110001001110001010001100101101010011010000101101111011100010000001011110001111110010010001100100110100011101001000001101110010100110001001010101 || !detection)
      failures = failures+1;

    received <= 542'b01000110001100001111011111100000111110101111001111100010001110001010100101101101001110010000011100000110100101110110001111010010110000110000001101011110000111011011000110101001010100100001100110111011011111100000010001001110000100101110111011110010101111111010010111011011111000011110100010100101001011011111010011110111001001010100100011100010110010010111111000110110111000111000101001111101101011000011111100001100010010001111111000111011101010110111110001110000001101011011011111101011001111011100100001001001101000001101100000100011011011;
    #1;
    if (message != 512'b01000110001100001111011111100000111110101111001111100010001110001010100101101101001110010000011100000110100101110110001111010010110000110000001101011110000111011011000110101001010100100001100110111011011111100000010001001110000100101110111011110010101111111010010111011011111000011110100010100101001011011111010011110111001001010100100011100010110010010111111000110110111000111000101001111101101011000011111100001100010010001111111000111011101010110111110001110000001101011011011111101011001111011100100001000001 || !detection)
      failures = failures+1;

    received <= 542'b01000111101010110110111100010000010011101100010100110100010111000001010011100001101001000000110101010010101001111000100110100110101101001110101010000110010101001001011110111000111101110110001101111001101100000011111011001000100011001011001011010100110000110101000001100100010001111110110101100010101111101100111101100011110111111001010110011111001101100000010100101001010101111011101100000101001110101101011110110010000110101110011011100011100110001101110101110111010010100010001001010000011101010000101100111000110010101101001111100001110100;
    #1;
    if (message != 512'b01000111101010110110111100010000010011101100010100110100010111000001010011100001101001000000110101010010101001111000100110100110101101001110101010000110010101001001011110111000111101110110001101111001101100000011111011001000100011001011001011010100110000110101000001100100010001111110110101100010101111101100111101100011110111111001010110011111001101100000010100101001010101111011101100000101011110101101011110110010000110101110011011100011100110001101110101110111010010100010001001010000011101010000101100111000 || !detection)
      failures = failures+1;

    received <= 542'b10111110011101110101000110010000101001000110011000001011111110000001101111110101101100011101001001100000100101001011010011110110010000001110101001100000010001001100000011111000100011010011000000111100000111100000100111111000111010110001111111111010000101111001001001011001010111101010110000000011100010000011001110110001010110011111100001100101011001011010001010000111010111111011110001000100110001010111111000110001011000110111111100011001101011000101010100001010001111110011111010011100000010011111010000100010110100111101000111010001101100;
    #1;
    if (message != 512'b10111110011101110101000110010000101001000110011000001011111110000001001111110101101100011101001001100000100101001011010011110110010000001110101001100000010001001100000011111000100011010011000000111100000111100000100111111000111010110001111111111010000101111001001001011001010111101010110000000011100010000011001110110001010110011111100001100101011001011010001010000111010111111011110001000100110001010111111000110001011000110111111100011001101011000101010100001010001111110011111010011100000010011111010000100010 || !detection)
      failures = failures+1;

    received <= 542'b11011001010000101101011110100000000111011101100111000010101001101101010000001100010000010110100000111011010011011101000101010010001011011010101001011111111101111110100000010010100111111011011101100000011111110100110101011010010001001010110011110111001011001000001010100000000011001111001100111000000000100101001001001011011010110110001110100100001111101111001101111001100011011110101001010101010001000101010100100111001101111010011000101111010001001101001100000111110101111010001110000100001100011100000100000111011110101001110100011010111101;
    #1;
    if (message != 512'b11011001010000101101011110100000000111011101100111000010101001101101010000001100010000010110100000111011010011011101000101010010001011011010101001011111111101111110100000010010100111111011011101100000011111110100110101011010010001001010110011110111001011001000001010100000000011001111001100111000000000100101001001001011011010110110001110100100001111101111001101111001100011011110101001010101010001000101010100100111001101111010011000101111010101001101001100000111110101111010001110000100001100011100000100000111 || !detection)
      failures = failures+1;

    received <= 542'b10001101111001000100101010001010101110110011101101111101100011000000100101011001000110100101111101011110110110110000001100110011100110110110011100100111010111001100101100011001001110111100000101111000111101001111000001010100010100110011110100101111111010110001010000111100101111001001001011110010001011111101001111011011101100101110110011110000100001110010111111000101010110001101001000010010011100100010100110001101100111001010110100001011011010111100010010001100011011010011111000001100110100001100110110001100001100111000111100000100101010;
    #1;
    if (message != 512'b10001101111001000100101010001010101110110011101101111101100011000000100101011001000110100101111101011110110110110000001100110011100110110110011100100111010111001100101100011001001110111100000101111000111101001111000001010100010100110011110100101111111010110001010000111100101111001001001011110010001011111101001111011011101100101110110011110000100011110010111111000101010110001101001000010010011100100010100110001101100111001010110100001011011010111100010010001100011011010011111000001100110100001100110110001100 || !detection)
      failures = failures+1;

    received <= 542'b00101110111101101100100010111101111100011011100110010111100001011110101001011111100010011000000001010001000100101010101101111100100000110101100010100011101000111110000100010001011110101101001110100101100001001110010011101111010010000101000100000101101000010111000011010111111010000110100001111011110010001001101001110101101110100010111000100011001001111011110100100001100011100010001110010101100001110110100010101010011001100010110011110000010100100010101010100101111000100110101100111011100111111001011101001111111000110100010110101011000011;
    #1;
    if (message != 512'b00101110111101101100100010111101111100011011100110010111100001011110101001011111100010011000000001010001000100101010101101111100100000110101100010100011101000111110000100010001011110101101001110100101100001001110010011101111010010000101000100000101101000010111000011010111111010000110100001111011110010001001101001110101101110100010111000100011001001111011110100100001100011100010001110010101100001110110100010101010011001100010110011110000010100100010101010100101111000100110101100111011100111111001011101001111 || !detection)
      failures = failures+1;

    received <= 542'b10010110101010011100011011101011111010011101101100010101100101000001010101110001001100101010011110010100101101100110100000101101110000100010011001011100000100111111010010010100000001011001010111100001001110001100111000011100000010111111100101101011010000110011001000101101000110110110011010011011000110111000101000010000100010101000001000011110101111010001000101000010000101010000001101110111010000000110001001110001100001011001111011001011110000101110101000011100000111100010110010101001010110001001100011111100100111101110000001000001111001;
    #1;
    if (message != 512'b10010110101010011100011011101011111010011101101100010101100101000001010101110001001100101010011110010100101101100110100000101101110000100010011001011100000100111111010010010100000001011001010111100001001110001100111000011100000010111111100101101011010000110011001000101101000110110110011010011011000110111000101000010000100010101000001000011110101111010001000101000010000101010000001101110111010000000110001001110001100001011001111011001011110000101010101000011100000111100010110010101001010110001001100011111100 || !detection)
      failures = failures+1;

    received <= 542'b01100001110100001100101101111111001100010101001111011010101110011001001111110111010010100111110001011101011011010011110001110100100110000011110010010101100110101110000100011010111101110000100000100101110001000111000000110000000011110011000111011001000010001111101100001000001100110001101011100001100110111100111101000101000010000010110010100100110110011101011101000011010110010001000001010110010101000000101111110110111110100010101001011000111100011001110000110100111101111010000010100000111111111111001001100110001010100010000100011011001110;
    #1;
    if (message != 512'b01100001110100001100101101111111001110010101001111011010101110011001001111110111010010100111110001011101011011010011110001110100100110000011110010010101100110101110000100011010111101110000100000100101110001000111000000110000000011110011000111011001000010001111101100001000001100110001101011100001100110111100111101000101000010000010110010100100110110011101011101000011010110010001000001010110010101000000101111110110111110100010101001011000111100011001110000110100111101111010000010100000111111111111001001100110 || !detection)
      failures = failures+1;

    received <= 542'b11001110101111010000011000011010110010001001100101100000011010010100111110111111001110001010110011110100110101001101010100111110111001111010011010011010110110001100001100100000111110101010011111101001110001001001001011000000110010101000100100011111011000000100010010110010001100011001110110011001001011010111101101101110011001110110110011100101101101101010011011010101111010001000010011001001010101100011001001011111000111011010001010010000100110100011111000010011110001011111000001100000101111010000010111100111100110111110000101101111111001;
    #1;
    if (message != 512'b11001110101111010000011000011010110010001001100101100000011010010100111110111111001110001010110011110100110101001101010100111110111001111010011010011010110110001100001100100000111110101010011111101001110001001001001011000000110010101000100100011111011000000100010010110010001100011001110110011001001011010111101101101110011001110100110011100101101101101010011011010101111010001000010011001001010101100011001001011111000111011010001010010000100110100011111000010011110001011111000001100000101111010000010111100111 || !detection)
      failures = failures+1;

    received <= 542'b01111100000011000011101101001000000111010110011010001110100000100101101010000110111100111100001011010011010001110011110101011111101101000111010011101110000111110100111011000111011110111111011111000100110111000011111011011011011010111101111001010010011001000101011010101010000111001101001001101011011010110101011010110101101001011011000100101101110010001111000101001111110011000010100001001111100110011111111010001101111001011001001010010100100010110101110010011010110000000110101010010000110000110100110100100011011100110010110111001111001000;
    #1;
    if (message != 512'b01111100000011000011101101001000000111010110011010001110100000100101101010000110111100111100001011010011010001110011110101011111101101000111010011101110000111110100111010000111011110111111011111000100110111000011111011011011011010111101111001010010011001000101011010101010000111001101001001101011011010110101011010110101101001011011000100101101110010001111000101001111110011000010100001001111100110011111111010001101111001011001001010010100100010110101110010011010110000000110101010010000110000110100110100100011 || !detection)
      failures = failures+1;

    received <= 542'b01110101001111110011100111111110000110011111111101100010110001011011100100010110010010111101100111100111001010110101110110011011111111100010001111011111110110000001011110100011100001110100000000100110111111001111111010100011111001000111000111101001111011111010110110100010111100000000010110011101001001110011011000001101011001110101111000101001111010011110011111111001110101110100010010011111100011100000001101011011000111101011001101001000001000011101101011111100111101000101001111101001000111000001111101101100101000101011000011011110011110;
    #1;
    if (message != 512'b01110101001111110011100111111110000110011111111101100010110001011011100100010110010010111101100111100111001010110101110110011011111111100010001111011111110110000001011110100011100001110100000000100110111111001111111010100011111001000111000111101001111011111010110110100010111100000100010110011101001001110011011000001101011001110101111000101001111010011110011111111001110101110100010010011111100011100000001101011011000111101011001101001000001000011101101011111100111101000101001111101001000111000001111101101100 || !detection)
      failures = failures+1;

    received <= 542'b11101100111100101000101111110011110110000001110110001010111010100000110000101101010000111101100001110001110110110010101111110010000101011011111100010100110010010011101010010101110001001011000111111110000001001000010111000100111110111011011010000011111100111111001101001110110011010000011100101111010011101001000101111010010111111101011011100110100100001001100100011101111000101000100010111100110000100110000011100101111010010000001111010110111110001010111111010100111011101100110110000001010100000010000101001010110010101100111010111100001100;
    #1;
    if (message != 512'b11101100111100101000101111110011110110000001110110001010111010100000110000101101010000111101100001110001110110110010101111110010000101011011111100010100110010010011101010010101110001001011000111111110000001001000010011000100111110111011011010000001111100111111001101001110110011010000011100101111010011101001000101111010010111111101011011100110100100001001100100011101111000101000100010111100110000100110000011100101111010010000001111010110111110001010111111010100111011101100110110000001010100000010000101001010 || !detection)
      failures = failures+1;

    received <= 542'b00001101111001111111001010100101000101111001001110111010000011010100111110000010001011110010111000010110010000111011010101100111100101101010101110101001110000111111000101110011000111111001101001100111110110100111001111110101101100001001010110000001000001100011011111110101000000101101100011001100101100010010010001010111001000101101101111000101110110101011110101110001111101010010010100000100011110111011101011000000010001110111101001001101101111101101011101100101101100110111101111111001110101111100101111110101001010000111001110010101110111;
    #1;
    if (message != 512'b00001101111001111111001010100101000101111001001110111010000011010100111110000010001011110010111000010110010000111011010101100111100101101010101110101001110000111111000101110011000111111001101001100111110110100111001111110101101100001011010110000001000001100011011111110101000000101101100011001100101100010010010001010111001000001101101111000101110110101011110101110001111101010010010100000100011110111011101011000000010001110111101001001101101111101101011101100101101100110111101111111001110101111100101111110101 || !detection)
      failures = failures+1;

    received <= 542'b00001101110101000001101101000010000010011110100111001111000111100010110101011010100101011010111011011000011111000101110000010010101111110100101000000101010010011011101010000001100010010011011110010110111100011010011110001101100000011010000110111000110101000111010010110010001100111000000000111100101001011001110101101000111001101000111101101111101010000101110100101110101011101001011000001110101010010111101100011000001011110100000011111010010010110100101101100101000011010100110010010101100000010101110001011101001101000011010101001001110001;
    #1;
    if (message != 512'b00001101110101000001101101000010000010011110100111001111000111100010110101011010100101011010111011011000011111000101110000010010111111110100101000000101010010011011101010000001100010010011011110010110111100011010011110001101100000111010000110111000110101000111010010110010001100111000000000111100101001011001110101101000111001101000111101101111101010000101110100101110101011101001011000001110101010010111101100011000001011110100000011111010010010110100101101100101000011010100110010010101100000010101110001011101 || !detection)
      failures = failures+1;

    received <= 542'b10000111000100100101110010011100010110101001111001001111011110011010001011011000001001011000100110010010110000001101001010000100111100101100010100101101111111101101111111010011111011001001011000100101111000100000011110011000001011000111101010001101000011001011010100010000010011011011100011111100001011101010001100100010011000001101110110101010010011010000101011011011111011111011001000111011010110000111111011001111110001111001000010011100111111111011100010011101110111010000111111111000110000111110001011100111100111000111110110011100101010;
    #1;
    if (message != 512'b10000111000100100101110010011100010110101001111001001111011110011010001011011000001001011000100110010010110000001101001010000100111100101100010100101101111111101101111111010011111011001001011000100101111000100000011110011000001011000111101010001101000011001011010100010000010011011011100011111100001011101010001100100010011000001101110110111010010011010000101011011011110011111011001000111011010110000111111011001111110001111001000010011100111111111011100010011101110111010000111111111000110000111110001011100111 || !detection)
      failures = failures+1;

    received <= 542'b11000101011110101101001011001100100110001111000010001110101010101110011111001111111111011011101110011100001010011010001001000100001010100100101011000101111000011000000001100000000001111001011111010101000001011010000110010010010011010001001101110100110000010010001011001000001110000010100011110111010101010011000000010001001110110011000100011011010111001100010010010011101100000111010101100000100111001110011011110110110010011001101001001111101000101011110011110010110110000001010101101111000100000011111100010110100111110100111100111000111100;
    #1;
    if (message != 512'b11000101011110101101001011001100100110001111000010001110101010101110011111001111111111111011101110011100001010011010001001000100001010100100101011000101111000011000000001100000000001111001011111010101000001011010000110010010010011010001001101110100110000010010001011001000001110000010100011110111010101010011000000010001001110110011000100011011010111001100010010010011101100000111010101100000100111001110011011110110110010011001101001001111101000101011110011110010110110000001010101101111000100000011111110010110 || !detection)
      failures = failures+1;

    received <= 542'b01001010011101000010011001100100100001001001110101111111001011010011000001011101110011011111111110111001101000111001111100000010101001000101001100111100110000111001010010110011111101010001110101011111001111001101111010100001000001011010111000000010100110010010010011001100101000101000100110000110101010111110000110111100111101111000001000010011000101001010011100011011101000101110110000100110111101100101100000101011000100010100110000010010111110101110100011110001000010111101100011010100010111100000110000100100001001000010101011010011000011;
    #1;
    if (message != 512'b01001010011101000010011001100100100001001001110101111111001011010011000001011101110011011111111110111001101000111001111100000010101001000101001100111100110000111001010010110011111101010001110101011111001111001101111010100001000001011010111000000010100110010010010011001100101000101000100110000110101010111110000110111100111101111000001000010011000101001010011100011011101000100110110000100110111101100001100000101011000100010100110000010010111110101110100011110001000010111101100011010100010111100000110000100100 || !detection)
      failures = failures+1;

    received <= 542'b01000111101000101110000000011110101011100000111000111000001111100111111110000000010100101000111010001000011111001000001001000011101110100111100100111010111000111001011100100110010000010000111000100110100011001111100011100001010011001111111011010111001110101101100001010001111111000101101010011011010100110100111111111111011111011001101110101100010100110101100111011000110110111001000010110100110100111110010000100111110110000101111110001100010101010010010100010001001110101111111001000111110110100000101110011111001011110101011011000011001010;
    #1;
    if (message != 512'b01000111101000101110000000011110101011100000111000111000001111100111111100000000010100101000111010001000011111001000001001000011101110100111100100111010111000111001011100100110010000010000111000100110100011001111100011100001010011001111111011010111001110101101100001010001111111000101101010011011010100110100111111111111011111011001101110101100010100110101101111011000110110111001000010110100110100111110010000100111110110000101111110001100010101010010010100010001001110101111111001000111110110100000101110011111 || !detection)
      failures = failures+1;

    received <= 542'b10110011000101000100101101101110001100100111111101101101101000101001110100110110010101111000101101010010001110101010111100001111101010001001100101001111010001111011111011111101001001110010101101111110010010100011001010101110011101011000110111110110000101111011110110101011111111000000110001000111001000010101110000111011101101001100010101110001001000001011100011100111010000010000100110111010101100101111011101101011000000001110100011100100101100000111001110111110011001110110110111100001011010100001011001110110100111101111111010100000000111;
    #1;
    if (message != 512'b10110011000101000100101101101110001100100111111101101101101000101001110100110110010101111001101101010010001110101010111100001111101010001001100101001111010001111011111011111101001001110010101101111110010010100011001010101110011101011000110111110110000101111011110110101011111111000000110001000111001000010101110000111011101101001100010101110000001000001011100011100111010000010000100110111010101100101111011101101011000000001110100011100100101100000111001110111110011001110110110111100001011010100001011001110110 || !detection)
      failures = failures+1;

    received <= 542'b00000100001100011010010101111001010011111001011110010100011000000111011001000001100110010010000011010010000000011001011000011001111100110100001010000001011001000100001110101011101111010011010011101110011110011010010001001111001001101001100110010011110111010001011001010010000001111010101110011101001101101001000110010001000110011001100000111100001001000011010001100010000001010100010010010111001000110011000110100011011000000101010000010011011111101010001100110000011110011110001110000000110000110101100100011001101110111111110101001100111001;
    #1;
    if (message != 512'b00000100001100011010010101111001010011111001011110010100011000000111011001000001100110010010000011010010000000011001011000011001111100110100001010000001011001001100001110101011111111010011010011101110011110011010010001001111001001101001100110010011110111010001011001010010000001111010101110011101001101101001000110010001000110011001100000111100001001000011010001100010000001010100010010010111001000110011000110100011011000000101010000010011011111101010001100110000011110011110001110000000110000110101100100011001 || !detection)
      failures = failures+1;

    received <= 542'b11000101100111110010011011001010111111011011001001011001000110011011100100111101110010110111010011010000010001101100010000011011001000111110101000000001100101001101000110001101001011000001011001101110100101010000100011000111010100001011010011010111001111010101100110111001110111011011011100110101001010110100100100010101110011010001000101011100100011111000111110111100001010100100111000000010111000110110101011000000101000001101110000110000101101001101100010111111101110100100100101011010011010010011110111010111110010001001110111100010001010;
    #1;
    if (message != 512'b11000101100111110010011011001010111111011011001001011001000110011011100100111101110010110111010011010000010001101100010000011011001000111110101000000001100101001101000110001101001011000001011001101110100101010000100011000101010100001011010011010111001111010101100110111001110111011011011100110101001010110100100100010101110011010001000101011100100011111000111110111100001010100100111000000010111000110110101011000000101000001101110000110000101101001101100010111111101110100100100101011010011010110011110111010111 || !detection)
      failures = failures+1;

    received <= 542'b00110000110111110001101111110000101101110001110110010100111010010101000111111101011000001010010011100111111111100000101101010110010011000011001110101100111000011110010000100100000111100001001000010101010011000100010010010101101001110100110101111011000101111011101001111010110101000001000101110011100101110000110101001100010100000110111110100010110010011110100001111000111010110111101110111000111100000100101101110111100001111110001001000000100111101000011010001101000011001010111110111010010011011111101000100101110100010010111000110011011011;
    #1;
    if (message != 512'b00110000110111110001101111110000101101110001110110010100111010010101000111111101011000001010010011100111111111100000101101010110010011000011001110101100111000011110010000100100000111100001001000010101010011001100010010010101101001110100110101111011000101111011101001111010110101000001000101110011100101110000110101001100010100000110111110100010110010011110100001111000111010110111101110111000111100000100101101110111100001111110001101000000100111101000011010001101000011001010111110111010010011011111101000100101 || !detection)
      failures = failures+1;

    received <= 542'b01000100100010000011000101000011000110111101000111001000110101111011010011001000010001110110110000101011110100100101000010111001010000110001001101110011011010111101101011011110011101111101110111011100000101111000010100010001101011011100111000111010101101010110111000011100001010101000011110010010001100101100010100101100110010000001111100101111011110101000111101010110000100011011011110110111111101100101111101101001110011101110000101101000011111111000011001100011000110010111011110001011000110011001110100111100010101111010110100111101011110;
    #1;
    if (message != 512'b01000100100010000011000101000011000110101101000111001000110101111011010011001000010001110110110000101011110100100101000010111001010000110001001101110011011010111101101011011110011101111101110111011100000101111000010100010001101011011101111000111010101101010110111000011100001010101000011110010010001100101100010100101100110010000001111100101111011110101000111101010110000100011011011110110111111101100101111101101001110011101110000101101000011111111000011001100011000110010111011110001011000110011001110100111100 || !detection)
      failures = failures+1;

    received <= 542'b10000101101000101101110011011110111011010001011001010100010101010100001011100111011011101100101010001110100101110011111011111011011010001011001010011011110010101110011011110001010100000100101111101101101010101100100110011111111101110001110111011001100101111100111100111111101011011100011001110011110111110001110111101001000001011000101001010100010100111010001110010011110000111011011001000010011111001011010101111100110001011101001001110101111011111000000001001111001000011110110101011011010111010110100010100100000001101000101010100011000001;
    #1;
    if (message != 512'b10000101101000001101110011011110111011010001011001010100010101010100001011100111011011101100101010001110100101110011111011111011011010001011001010011011110010101110011011110001010100000100101111101101101010101100100110011111111101110001110111011001100101111100111100111111101011011100011001110011110111110001110111101001000001011000101001010100010100111010001110010011110000111011011001000010011111011011010101111100110001011101001001110101111011111000000001001111001000011110110101011011010111010110100010100100 || !detection)
      failures = failures+1;

    received <= 542'b00001001010000101111000101100010100001111100001110111111111100011011100010001110010101101000000001000110010111111111110101011111011100001110100010010110001100101001011111100101000101101100100011101111000001000010010110000100111110110011011010011000111000001000001100100111110001111001101011111010010101011010011100101010010011000010111110001110001111001000110111110110110111010101010101001111111000101011010110111001111100111000111110001110100000000101000100010101000101101000100100100000011010010000100110010101011100111001011011001010000110;
    #1;
    if (message != 512'b00001001010000101111000101100010100001111100001110111111111100011011100010001110010101101000000001000110010111111111110101011111011100001110100010010110001100101001011111100101000001101100100011101111000001000010010110000100111110110011011010011000111000001000001100100111110001111001101011111010010101011010011100101010010011000010111110001110001111001000110111110110100111010101010101001111111000101011010110111001111100111000111110001110100000000101000100010101000101101000100100100000011010010000100110010101 || !detection)
      failures = failures+1;

    received <= 542'b01100110100010111010010010010010100010110001100001110001000010101100010100010000010101111000100000010001111000011111100000011000011010001101011000000110111000000100011100001001010101011110011011110001000101101010011110100000001100110001011000011011100010001101011001110111000111001101111101010111000110100100010111110011010000011000001100110001100110001110101010111110101101101010011111001000101101010010010111111010100010010001101100101100100101101011101010001011101101110001110110100001001110100010110111111100101101101001010010011101010011;
    #1;
    if (message != 512'b01100110100010111010010010010010100010110001100001110001000010101100010100010000010101111000100000010001111000011111000000011000011010001101011000000110111000000100011100001001010100011110011011110001000101101010011110100000001100110001011000011011100010001101011001110111000111001101111101010111000110100100010111110011010000011000001100110001100110001110101010111110101101101010011111001000101101010010010111111010100010010001101100101100100101101011101010001011101101110001110110100001001110100010110111111100 || !detection)
      failures = failures+1;

    received <= 542'b10010011000000100111001101100110111110000101100110001111011011010011010101001111101010010101100111011000111111000011000100001011110010111000010111001011010011000011101011001110111101010100100011010011100001100001101001101101011110001001011010001100101111011110100110000110000110001001011010101011011001000110001101110001101011011010101010010100110100101110111010110001000001101010101101111111101100110010100010010000100101110111111010100000001011010101001100000011100000101100111000011100111011011110100111001001110011101001101101000001010101;
    #1;
    if (message != 512'b10010011000000100111001101100110111110000101100110001111011011010011010101001111101010010101100111011000111111000011000100001011110010111000010111001011010011000011101011001110111101010100100011010011100001100001101001101101011110001001011010001100101111011110100110000110000110001001011010101011011001000110001101110001101011011010100010010100110100101110111011110001000001101010101101111111101100110010100010010000100101110111111010100000001011010101001100000011100000101100111000011100111011011110100111001001 || !detection)
      failures = failures+1;

    received <= 542'b00110000101010100000110100111100110001001010101100010101110010111110011010100101001000010010111011101010000010011100111010000111100001000101011010111010010011111001101001101010111101110010001001000110000010000110001000010010101010100000001111100100100101110101010010011011110010111110000011110111111100000000010000000101001101110001011001110000001101011011110001111001001110000010100011001011000101010010111000100101001100100010110100011100000110000010110101000110110000101010000011110000001100101000011000001011011100111001000001000101010100;
    #1;
    if (message != 512'b00110000101010100000110100111100110001001010101100010101110010111110011010100111001000010010111011101010000010011100111010000111100001000101011010111010010011111001101001101010111101110010001001000110000010000110001000010010101010100000001111100100100101110101010010011011110010111110000011100111111100000000010000000101001101110001011001110000001101011011110001111001001110000010100011001011000101010010111000100101001100100010110100011100000110000010110101000110110000101010000011110000001100101000011000001011 || !detection)
      failures = failures+1;

    received <= 542'b11011001100010011110001001001110110100001010110000110100100001011001011010111010010110001110110010010111011110000110100010000001100100011111001110111100110000111011100010010110011101100100100000010011101001110010010110001100100010111010110011101110110001011111100100110101010101001000001100100011100100001000100101101000100000000111100000011010000011100111010110110100100010101110010110111011101100000010101010011101101001100111101011100110010011000101000111011101100111011000011001110111001101000100110110001011110111001101000100001100001100;
    #1;
    if (message != 512'b11011001100010011110001001001110110100001010110000110100100001011001011010111010010110001110110010010111011110000110100010000001100100011111001110111100110000101011100010010110011101100100100000010011101001110010010110001100100010111010110011101110110001011111100100110101010101001000001100100011100100001000100101101000100000000111100000010010000011100111010110110100100010101110010110111011101100000010101010011101101001100111101011100110010011000101000111011101100111011000011001110111001101000100110110001011 || !detection)
      failures = failures+1;

    received <= 542'b11110110011010101111000110010000000000000110110010010010110011010110101010010111111011000011111001011011010001100110110110111101111100000100001010011100100001110110000111111101100010100011111111010110101010101110000111000011010111110010010010111010100001110110100010101001011011011010110010101001010110110101010011110010001011001110100111010000110010011000011010101101110100001101110101101001110110111110100001000110100011110011011100110000001001011001110000100011011010001000111010110110010111010111111101000100100011110000110001111110101111;
    #1;
    if (message != 512'b11110110011010101111000110010000000000000110110010010010110011010110101010010111111011000011111001011011010001100110110110111101111100000100001010011100100001110110000111111101100010100011111111010110101010101110000111000011010111110010011010111010100001110110100010101001011011011010110010101001010110110101010011110010001011001110100111010000110010011000011010101101110100001101110101101001110110111110100001000110100011110011011100110000001001011011110000100011011010001000111010110110010111010111111101000100 || !detection)
      failures = failures+1;

    received <= 542'b11110101110011111010101110111001111001001010000101011101001001100101000000010110011101100100100011001100100010111111001000000101100111100001011001011001010110110001010010111111111101111011111100101001000010010111100001000110011000011000101100000001110111110010010001101000010001100101011101111101110110101000010011010011111100001010000001000010110000010110111100011001011111011010000111110111100011100101000000000001000010101110101001010010111011000101100110101111000111110100100001010000001100111100100000000010001001110010100111011110101010;
    #1;
    if (message != 512'b11110101110011111010101110111001111001001010000101011101001001100101000000010110011101100100100011001100100010111111001000000101100111100001011001011001010110110001010010111111111101111111111100101001000010010111100001000110011000011000101100000001110111110010010001101000010001100101011101111101110110101000010011000011111100001010000001000010110000010110111100011001011111011010000111110111100011100101000000000001000010101110101001010010111011000101100110101111000111110100100001010000001100111100100000000010 || !detection)
      failures = failures+1;

    received <= 542'b11000001001010010101101110111011001111110111010000010111000100110011010111000011010110100111110011010101110110001001010010100110010011101010100001001111010000101011111010010100010111001001000110100111011010010111110001110000101010110010001001101001010010110111100110100001011000111000011001001010010011111010011011000101101000100100010110000000111001100110001111111000101100011100010111110110001001110011001100110010000011101111111011011011000001101111001011010010011000000001111111011101010111000000010110010010111101101010000100110101001111;
    #1;
    if (message != 512'b11000001001010010101101110111011001110110111010000010111000100110011010111000011010110100111110011010101110110001001010010100110010011101010100001001111010000101011111010010100010111001001000110100111011011010111110001110000101010110010001001101001010010110111100110100001011000111000011001001010010011111010011011000101101000100100010110000000111001100110001111111000101100011100010111110110001001110011001100110010000011101111111011011011000001101111001011010010011000000101111111011101010111000000010110010010 || !detection)
      failures = failures+1;

    received <= 542'b01110100001101001001000000010001111000110111010100000000001010010010110111001110011001111010011010011000101011000101110111111100001111100001100010111111000110000010010110110100011001101110010101101011111101110111101101101010000100111010101101011100001100101100110110011011100011011110011110100011100001011101101100010001000010000101101001101001101010100101000000010001100101100110110111100100110001100101100001000001111010000100110101111100111011100100011010111010000101000010111011111100111100001010111110110010000011111000101100111010010011;
    #1;
    if (message != 512'b01110100001101001001000000010001110000110111010100000000001010010010110111001110011001111010011010010000101011000101110111111100001111100001100010111111000110000010010110110100011001101110010101101011111101110111101101101010000100111010101101011100001100101100110110011011100011011110011110100011100001011101101100010001000010000101101001101001101010100101000000010001100101100110110111100100110001100101100001000001110010000100110101111100111011100100011010111010000101000010111011111100111100001010111110110010 || !detection)
      failures = failures+1;

    received <= 542'b11111011000001000001110101000010011110001010101101000110011010110001100000011001010111100010010111100011011011010000101101100100011001101000101000100010010101001111001101110100011101111111011111100100001010000000100100010001101100111010011010011110110001001000010000001111111011010100111101111001000100000001100010101011111100110000101101100001110000001110000011111001101111011011000110101110000111100111101010101100101100001000110001110000011000001110100000100100101010111100111111101111000011111101110110100010011100110111110111111011110100;
    #1;
    if (message != 512'b11111011000001000001110101000010011110001010101101000110011010110001100000011001010111100010010111100011011011010000101101100100011001101000101000100010010101001111001101110100011101111111011111100100001010000000100000010001101100111010011010011110110001001000010000001111111011010100111101111001000100000001100010101011111100110000101101100001110000001110000011111001101111011011000110101000000111100111101010101100101100001000110001110000011000001110100000100100101010111100111111101111000011111101110110100010 || !detection)
      failures = failures+1;

    received <= 542'b11010110100000001110110010011101101011011000001100100000010001010011100110110101101111100001111100101100011010110011111010011110010101101101101110111010111101000010001011101001101100110110110011111000010010110001111110011011100111000010010101011000010001111011110010101001001101010011111010001110111110111000011110111110100101110110101110010101111111010011000011010010010010010011110100100110100101000011000011000010011101101100100111100011010001101110001100011101000100101000100110101010100111110010010101011101010001010101111010000111001000;
    #1;
    if (message != 512'b11010110100000001110110010011101101011011000001100100000010001010011100110110101101111100001111100101100011010110011111010011110000101101101101110111010111101000010001011101001001100110110110011111000010010110001111110011011100111000010010101011000010001101011110010101001001101010011111010001110111110111000011110111110100101110110101110010101111111010011000011010010010010010011110100100110100101000011000011000010011101101100100111100011010001101110001100011101000100101000100110101010100111110010010101011101 || !detection)
      failures = failures+1;

    received <= 542'b00100110101101010000000101101000100010011101000000010111001111011100000010101011111011001100000001110000011100011001110110001101101110111001001010000100100001001111100000111010010000100101011010101110100010111010001111100011101011010101100101000001011010101001110010010111011011010011110001110010101100001011100010001000110100101101000011000011101101010011111011011101101000111111100001100000000111001011010010110111000011101110100011011000100101110110100001100001111110000011101001100011000100011100010000010111111010111011000100101000111000;
    #1;
    if (message != 512'b00100110101101010000000101101000100010011101000000010111001111011100000010101011111011001100000001110000011100011001110110001101101110111001011010000100100001001111100000111010010000100101011010101110100000111010001111100011101011010101100101000001011010101001110010010111011011010011110001110010101100001011100010001000110100101101000011000011101101010011111011011101101000111111100001100000000111001011010010110111000011101110100011011000100101110110100001100001111110000011101001100011000100011100010000010111 || !detection)
      failures = failures+1;

    received <= 542'b11101111001011110001110010110100100010101010100101101111110101011001100100111000101111100011001010100101010100110010010101010111010001111001110100010110011001010000001100010000111110011100010110000010011000010001011100101010100001011001111101011111001001110111011101011101010101111111100111001011100010011001111110010001011111000000011000000010111100001110010001110110001010111010111011111000010001001110000101110101110011001011110111010010101101010111001100111100001010101010101101100100110001110101101011000101000111001111001010110100000101;
    #1;
    if (message != 512'b11101111001011110001110010110100100010101010100101101111110101011001100100111000101111100011001010100101010100110010010101010111010001111001110100010110011001010000001100010000111110011100010110000010011000010001011100101010100001011001111101011111001001110111001101011101010101111111100111001011100010011001111110010001011111000000011000000010111100001110010001110110001010111010111010111000010001001110000101110101110011001011110111010010101101010111001100111100001010101010101101100100110001110101101011000111 || !detection)
      failures = failures+1;

    received <= 542'b10100100100010110000000101100010011101100101010101000111001001011010001100011101111011010010010001100001111110000011000110001000100101110010110000011100011001000011110001101100101111001010011101010000011010111101100001101110111000100011000011011001001000000000101010100011110010010000110011011111011011011101010010010110100101000100011001011010001111010111110000110001000111101010000110010100111111011010101101010011001010111000000111001111110010001001111111011101001111110101011000010100101011111111011001110001000101111001011101111100001011;
    #1;
    if (message != 512'b10100100100010110000000101100010011101100101010101000111001001011010001100011101111011010010010001100001111110000011000110001000100101110010110000011100011001000011110101101100101111001010011101010000011010111101100001101110111000100011000011011001001000000000101010100011110010010000110011011111011011011101010010010110100101000100011001011010001111010111110100110001000111101010000110010100111111011010101101010011001010111000000011001111110010001001111111011101001111110101011000010100101011111111011001110001 || !detection)
      failures = failures+1;

    received <= 542'b11100011010001100011010110000100001000110010001010111000101011110101001111110111000111001101010100010010011010101011111111001001110111001001000110000001000010001011110000000111100011111111001001010111100101100111110110100100001000000101001011001101000010001101110001000100010100011001111110100010011100000010100001011100101111000011011110010111101100100101110110101110111001000110000010001110001100000011001001010111110110010001100001111111010111000111011010110001011101110001101000001111010100110111011000011101100101011001100011111000111001;
    #1;
    if (message != 512'b11100011010001100011010110000100001000110010001010111000101011110101001111110111000111001101010100010010011010101011111111001001110111001000000110000001000010001011110000000111100011111111001001010111100101100111110110100100001000000101001011001101000010001101110001000100010100011001111110100010011100000010100001011100101111000011011110010110101100100101110110101110111011000110000010001110001100000011001001010111110110010001100001111111010111000111011010110001011101110001101000001111010100110111011000011101 || !detection)
      failures = failures+1;

    received <= 542'b11111111010010011000000100010110101100001000101010011111110101110001001011000010101011010010001101110111001000001011011000011011001100000001110001000110101001011001000001010000011010111101001110100111010100111100101001001010011110110001010111110000000000101000110011110001010111101101100001001100010101111111100011100011100011100100010101001000000010110010111001101101010101010011100011010011111101010100010011010010110101000110011001001100101110101010110110111100001001101001010110111001001100000011011001110011010110111001011100111100100111;
    #1;
    if (message != 512'b11111111010010011000000100010110101100001000101010011111110101110001001011000010101011010010001101110111001000001011111000011011001100000001110001000110101001011001000001010000011010111101001110100111010100111100101001001010011110110001010111110000000000101000110011110001010111101001100001001100010101111111100011100011100011100100010101001000000010110010111001101101010101010011100011010011111101010100010011010010110101000110011001001100101110101010110110111100001001101001010110111001001100000011011001110011 || !detection)
      failures = failures+1;

    received <= 542'b00001011001110110101010100011000000111011110001100111110100001001010110110100110110000101001001000000101001101110011110001100100010111000111111100101101110011110110101100011100100000010100010101111101111010001110000010010000110001101001110001000101010111101010110000001100010101110100101000100100110001101011110000110001001000011011010100100010011101001101100110101101101111111101010000000110111011100000011001101101000000011000000110100111110001001100101011101001001100000110011110000011001000001101001001011010010011001100011101111000011000;
    #1;
    if (message != 512'b01001011001110110101010100011000000111011110001100111110100001001010110110100110110000101001001000000101001101110011110001100100010111000111111100101101110011110110101100011100000000010100010101111101111010001110000010110000110001101001110001000101010111101010110000001100010101110100101000100100110001101011110000110001001000011011010100100010011101001101100110101101101111111101010000000110111011100000011001101101000000011000000110100111110001001100101011101001001100000110011110000011001000001101001001011010 || !detection)
      failures = failures+1;

    received <= 542'b01101111000001111010000000000111001111000010011111101000111011000111111010111100011001111100101011011000001001000011011011111010010111111111111110001101001100010110000100100010101111101110010000101111000111011110110101101000100110001111011100000110101111100010011101001100001101000011011010000100001111100011111001100100011011101011111011101100101000011100111111111000110011011101011111100000111001100101001110000001100000010101101101110010111011001110011110101011101011001001111110010010110011101011001011011101011010010111010101101101010001;
    #1;
    if (message != 512'b01101111000001111010000000000111001111000010011111101000111011000111111010111100011001111100101011011000001001000011011011111010010111111111111110001101001110010110000100100010101111101110010000101111000111011110110101101000100110001111011100000110101111100010011101001100001101000011011010000100001111100011111001100100011011101011111011101100101000011100111111111000110011011101011111100000111001100101001110000101100000010101101101110010111011001110011110101011101011001000111110010010110011101011001011011101 || !detection)
      failures = failures+1;

    received <= 542'b11101111110110010100100111010110010000001111011010000111100000111001000100100101101001111011101100010100001100101011010010100100101001010100101010111111101011010001110011100010011001010111111101001011101010000111101101001001000001011110101101011011110101100001010001001000011100110001010101110001001100110101111100001100110011110110110001100110110011011101100001111001100010001100100010100010011011100101101001101111100010101010010011001110111111111001100000101110010001100101001111001101011001011000111000001010010000111101110110001011010011;
    #1;
    if (message != 512'b11101111110110010100100111010110010000001111011010000111100000111001000100100101101001111011101100010100001100101011010010100100101001000100101010111111101011010001110011100010011001010111111101001011101010000111101101001001000001011110101101011011110101100001010001001000011100110001010101110001001100010101111100001100110011110110110001100110110001011101100001111001100010001100100010100010011011100101101001101111100010101010010011001110111111111001100000101110010001100101001111001101011001011000111000001010 || !detection)
      failures = failures+1;

    received <= 542'b01000101000100100101001100010111111110010011101001001111000110101111101000111101000000011001101011111000100100110111010100000011101111010101001000011111010101100011011110101011110001100001101000000110110010000110001011110011011001001001010110101001011000000100110111100000100011110001101101111000010000000011011000010000001111100111101111001110101001100110100101000000101100001111000110111011011001001001110110100001010100000011010000110111010101001110011100101100010101111011001010000001111101110011011101111001110110011100001101110001010100;
    #1;
    if (message != 512'b01000101000100100101001100010111111110010011101001001111000110101111101000111101000000011001101011111000100100110111010100000011101111010101001000011111010101100011011110101011110001100001101000000110110010000110001011110011011001001001010110101001011000000100110111100000100011110001101101111000010000000011011000010100001111100111101111001110101001101110100101000000101000001111000110111011011001001001110110100001010100000011010000110111010101001110011100101100010101111011001010000001111101110011011101111001 || !detection)
      failures = failures+1;

    received <= 542'b11101000110100100110000010100101001101100001101110000011011011000111101110000000011001100010111000110101110001010001011111100100010010110111111111000001101001000100100010100010010011110000111101110100000011100011100000110011100111010001010100010010011110000001100000101011110011000001011000110110010000111100111000000101100101010101011101000111000110110111100111000011001111000100000110100001001001111011100001000011010011010010011101100000000000111111001000111001101101001010100100100101111110010011010001110010000001101101101000111001101101;
    #1;
    if (message != 512'b11101000110100100110000010100101001101100001101110000011011011000111101110000000011001100010111000110101110001010001011111100100010010110111111111000001101001000100100010100010010011110000111101110100100011101011100000110011100111010001010110010010011110000001100000101011110011000001011000110110010000111100111000000101100101010101011101000111000110110111100111000011001111000100000110100001001001111011100001000011010011010010011101100000000000111111001000111001101101001010100100100101111110010011010001110010 || !detection)
      failures = failures+1;

    received <= 542'b00100100010111001101011111111001010111110110110111100101111101111011011010011100110100010111010100010111110010011111101101000110111010111101100100010001111101111110011111101001101101111101000001111011000101010010111110010001101001110100111100111010001011111111110100111111011001101001111000111110100110110110001010101101010111010101100101101111101011001101010010111001111000001000001010100100110100001101101000101001011001001111111011111000110100000001011001111111001011001101000000000000101100110111101010011100001001101001110110111010100111;
    #1;
    if (message != 512'b00100100010111001101011111111001010111110110110111100101111101111011011010011100110100010111010100010111110010011111101101000110111010111101100100010001111101111110011111101001101101111101000001111011000101010010111110010001101001110100111100011010001011111111110100111111011001101001111000111110100110110110001010101101010111010101100100101111100011001101010010111001111000001000001010100100110100001101101000101001011001001111111011111000110100000001011001111111001011001101000000000000101100110111101010011100 || !detection)
      failures = failures+1;

    received <= 542'b00010001001111110100110001101101110101101110000010110010110010101000000110000111010111011001010110011111110101110100111010110101001101000101000001010101100011001100110000000001000100011001011111111000010010111110000111100001000011010010100101111011101011001001011100011100011100100011101100010100000001110010001111101011010000011010000010101100000001111110000100011100101111111011111010010001111101011101000011101000001100001010101100100001010011011010111100101000111100000010010111100100000110011110101110010011111001000101010011010100000110;
    #1;
    if (message != 512'b00011001001111110100110001100101110101101110000010110010110010101000000110000111010111011001010110011111110101110100111010110101001101000101000001010101100011001100110000000001000100011001011111111000010010111110000111100001000011010010100101111011101011001001011100011100011100100011101100110100000001110010001111101011010000011010000010101100000001111110000100011100101111111011111010010001111101011101000011101000001100001010101100100001010011011010111100101000111100000010010111100100000110011110101110010011 || !detection)
      failures = failures+1;

    received <= 542'b00000011000010010010110010110011100111110010100100101010101010101000100111101000011011101111101100111101011110001110010111010000011101110111011101011011010100010001010000001011010000100010110101100100001000010000101011110111100000001010100010000111010101010111010001001111110001001010011000001101100000001101100101101101101000000000100110010010000110010100110000100111101000011100010100010011111100011100101000101011111010001101110000110001000001111100010011111000000100011111101110000010001010110111011000110010010101010101110110000110100100;
    #1;
    if (message != 512'b00000011000010010010110010110011100111110010100100101010101010101000100111101000011011101111101100111101011110001110010111010000011101110111011101011011010100010001010000001011010000100010110101100100001000010000101011110111100000001010100010000111010101010111010001001111110001001010001000001101100000001101100101101101101000000000100110010010000100010100110000100111101000011100010100010011111110011100101000101011111010001101110000110001000001111100010011111000000100011111101110000010001010110111011000110010 || !detection)
      failures = failures+1;

    received <= 542'b00111111011000011101110110010000101110111111011001100100001101011110110010011011000101110001010010110000011010100100000001101001011110100100000000110011000101101010001101100110110111111000011101111111000011100010100100010000010000000110000110011010110010000000011011111110000100101010011001100111000111100100011101100111001010010110001100001011101011100011010011111001010111000110100001111100011110000001100001111101010001101001110111110100111111000111001111100110000010011000110111110010111111001000000100100011110111001010101110000111110100;
    #1;
    if (message != 512'b00111111011000011101110110010000101110111111011001100100001101011110110010011011000101110001010010110000011010100100000001101001011110100100000000110011000101101010001101100110110111111000011101111111000011100010100100010000010000000110000110011010110010000000011011111110000100101010011001100111000111100100011101100111011010011110001100001011100011100011010011111001010111000110100001111100011110000001100001111101010001101001110111110100111111000111001111100110000010011000110111110010111111001000000100100011 || !detection)
      failures = failures+1;

    received <= 542'b11100001001000101010100110000111010111101011111110100010101110111101011110100101011010000100001100101100000001100010010001101010101001010001001101111001110110101101011001001110100001001001111111000101111001101111001100010110011010000011000111100001001010110010101010000100000001101100011011010000000110110000101011110110001000100001110110011110101100110001110101110010000101010011100110111010110001000111001011100001101010011101101000111000001001111111000010100000000111000111111000111011101100101000111000111110001100100101010001001010011100;
    #1;
    if (message != 512'b11100001001000101010100110000111010111101011111110100010101110111101011110100101011010000100001100101100000001100010010001101010101101010001001101111001110110101101011001001110110001001001111111000101111001101111001100010110011010000011000111100001001010110010101010000100000001101100011011010000000111110000101011110110001000100001110110011110101100110001110101110010000101010011100110111010110001000111001011100001101010011101101000111000001001111111000010100000000111000111111000111011101100101000111000111110 || !detection)
      failures = failures+1;

    received <= 542'b11111110110101010001010000100000000011001000111011110100101010001110101101111001110011110011110101010111011000110011011001010001110111000000111110001101000100010000110100101101010101000101110001100001110100101010011010101100010100000000100001010100101001010000110110100101000001101000101010000011001000100000101011101110110001011101111110000010011110110110100011110001010010000111000111110101100000101011000100000101100111001000111110100110010101100001010101101101101000001000101110000010000101100101000001011011110011101011110001001001001101;
    #1;
    if (message != 512'b11111110110101010001010000100000000011001000111011110100101010001110101101111001110011110011110101010111011000110011011001010001110111010000111110001101000100010000110100101101010101000101110001100001110100101010011010101100010100000000100001010100101001010000110110101101000001101000101010000011001000100000101011101110110001011101111110000010011110111110100011110001010010000111000111110101100000101011000100000101100111001000111110100110010101100001010101101101101000001000101110000010000101100101000001011011 || !detection)
      failures = failures+1;

    received <= 542'b01100110110011010000111010001010111110000010010110110000101101000010111011010010101010110111100101010010011011010011110010011101000000011001011001111000111111011111111000110001001100111000111000000110110010001110101000101111111000000011000110011100100010100110111110101101001111011011000110000000101011011001000000100100111111001000101010011101100011010111101000000111111101101100011010101011111000001001010110010101011101011011111001101000111010100111111100101100101011101011101111101111111111111001010100100100110111011110011110100100101110;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00110001110001011110001111100011000010100100010100000000110110011001101001100011111010000111011100010011101111111000111001001100011110010001100111100000001100111001000001000000011110110011100010100000001101111010101011111001000000111000100101010101110000111011111101011101010101111111001010001010111100101101101001101100011101010001111001110001100100100000011011000011001110111010000000100100010110001100101110001000011100110111111111111010101110000111101111010110111001101000111010111000000001110000001000100100111010111110100011011110111100;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00101000000101100000011011011011010111110101101010101001101101100110110101011101110111111100001011100011011100010110110111011101000101100100100001101000110000111001100110011111110011000010101101001110010101000011101110011110011110100010100011001010111101101111011001100010100100110010101111000110000001001100100000101110010101001111001011111100011010111110111100100111001001101100110110000000000001011011110000001100101000000011010001111110001000011110111100100100000111110011110111011010011100101100100101100000001110110110001010101110110011;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00011101110011101110010000000011110010100100001100000110110011110101110001000010101011100100110011100011000010111001010001000001011110100111100010111001100111000000010101100001000000000111000100111110011111010101001011111111010011101010000000111011111010000001000110101001110101111101010100000010001111110100011001110000101000101000100011010001010001110111100011111100010001010111011111110010110000010111011101000111100000001001111100000111111000011001110101101111111100011100100010100100010101101110010101001010010110010001111101100011000001;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b11011000111101101111000110100111101010110111100000001101011111110010110101001111000001000011110011111110101111001010001011010000011001101011110100001000110010100111110001011000001011010100101011000011000111101111100100011000011110111001110111110111011100100110000001100110100111110100000000011111111111010000001101100011101100001100010111011100010100111111100010100001000011101110111101011011010000001000011000101100101010100000110110000011111001101001010101001111000001000101111011001110001010100111111111111111110011111010110000011101101110;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00000110011100110010100010111001010001001101111011000100111110010000101110001101010000010110101101000111110100101000011001000111010000111111010100011011110110100001010110001001001010111110111100100101001001100111010001010110011001010011111000010101010111101000001110010100000111010100111010100101101011000101011001010000001101000010100010010111010011101100100101110011000001101000010011001100100100111101110011101101011000001001001010010001010100011110001000100101111101001011010001101110111011010010111000000111000000011110111110001101110010;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b11111000100101100101110111011101001001100011001010111000010001111110111010101111111000101101000101100010110111011011110110011010001110010111011110011100010101010110101111111100010100101000001100010110110111111100100101001110110100111000110010110011010011100100101010110011001111011010001110111111101100110101001101001010010000010011100001100100110100101100000010011111100100110111101001111100000101100011010101111101110110011110000010010001001000100110011111011101010000001001111110101100001010000100001110100111011010111010100000001100111011;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b01101000010110110001111011011011001100110101001101111000000011111100101101100011001011110101010000111110011110011100000110010011010100100101010110110000010111000011101010111100100101010101011101010101000111111001110100110001011110011001001111001010110010010111010011101001111100011000011111101000100100111010010101010101000100110100011110010010001101001110111101010101010111000100010000111010001101110100010001011110010000000010111001010001100001010101110011111010011101011010110011010001100000100100010100101001110001111111110010100111010010;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b01001010100011100001111011010111001011000110101111101000010001111010101111100011100111110001111111001011000101111111110010100100001111010010001001001110101110110101100111001101100111110000100101011110111011100111101000010010000101111000001010001011111010011001110111110000110011010110010110100100010110110100110101010111011100101101110100111011001010110110010001001110011101000001000000010110011000010111101101010111100001011000111100000011000000001000010111111000100110110100011000101100111101010111000001010111001011111001001011110101100101;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b01111100100001110111101110010110010101011101110110111001011110100111010110111100101111000101101000000001101001000011111010111011000011111101010110111000000010000001010010011011100101000111010110100101110011111110011110110010111001111111100110101100010100000010010101100110101110011011110110011011100111101101111000000100001111000011101111000110110101110000000010000101000011100101000010010100100001011100100000010000101001101011101101010011010101010001001010110100000011010111110000100011111100100101101101101000011101001011001000010010111000;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b10111010010100101111010100000111010110100111110011011100001010100100101011001100000000000101100110010101001101001000110100010000010011010111111010110010001011111111101001000110100000110001011000010011011001101001010000110010001011001110101000000011110010101001010100100011000000000010000110011001101110101000011110010110100100101111100001101110010100110010000010001111101000101000100000101011101010101101001011101010100001010111010100001100000010001001101100100111111100001011011010111001000111011111001101010001101110101101001101111000100010;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b01000000110101000100000010010111101101011000011001101001001001001001101000111010001110101001000110110110110111010000011011010001111100001010001111011100100000001000001011010001110000011011100000100010100000101001100101110011101011001010010101010000110100010101100010010101001101011011111000010100110000110001101000010011010010001000010100010110010010101111010000100111110000010100010010001101110111111101100100000011100111111101000000100101010010110001100011111000100010001100010111000011111101001110101100101001101110000101110100001100110001;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b10011001110001011111110010011101010011101100011101111111001111100111000111111001010011100111110111001110000000011111101010000111110100101000011111110100100000100111000001100110110000011011010001100111011011101000101011101010100100111001010111000110100001000011111011101000100101000000010100000101101001000001001000110111001110100000000100010101100100111110100101110100011000000011011010110110011001000101110100111100000011011111010101011010010001111101001010100010101001000110111010111111111011111010000100000001101101011110000110101100110110;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00101000011111000010011011000010111111100000110000100011001001011111101110100010100110101101110000100110010001000111000011110010011101101001010111000000001101110111011011011011101000111000100011011111010110110100011001000001110100101100101010100111010100110110000101111000100101011000011000100111010011110011010101001101010011001100000111001100100111010100010001011110000001110010100111111111000111010001100011110000111101011100100010000000101000110011100010001010100111111001000101111011111101011001100110011001101110100110110000001000101001;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00000011101011011110000001111001010101011010000101011001101110001101001101011010000101000101110111010001001001011110011101010101010101101001011100110111100100011010110010011000000100010101001101001001011111010101001101100111110000101110100110010011011100101101111001001110010010100000111010110100001111100100001010010111001101101011111001110001001011010010101100011111100011100000001000010010101101001010001001100101011101000100000000000001010111011111111001010010011110000101010111101110110010100000001101110101010010000001110001011110111110;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00001011000100001101100101111101011000000010111110001101100111101101011101001100001100110001011100001100101010111110100011010100111110000100000100111101000000010111001111101100010010111100111110000010011101001001000111011000101001110101001110101100000001010000010010010011111010000100011001000101101101001110101000010111100011101001100101101110001010101111001000111000010110011000000100101001000110000110110110101101000001100000111001000111000010110010011011110000111000000001110111010011100000000110001111101000010110001111100001011110110100;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b11001010111001100110001011000100101100000011010100101101100000100011010010110000101001010000101000101101111000110100100110001100010000100000100001110010111011110011010010110111010101100000010111011001111100000110000101010101101011001010000000011011110010110001011001110110101111010000101011010110001010100100100010000001111000110010010000010011000111101001011100001011111100011011101011001010000011011111011011111110011111110000110010011010101001001011001000100110000110100001011100101001000010000100000011111111110110100011000101011000001001;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b10010111010110011100101110110110001010010100000100110101100111010101111100000111010001001010110001101111011001101101111001010001011010000100111101010011110000010111101000110011100010011100111000110101001010111000100010010110010001100011010001101001000000001001010011000000011100111101110001001001001000111010111100110011101100111000111100101101100011110011011110101101111100101001000001111111100000010001100011010001101011001000001111010110001101001001010111110000000100000010101101010110100001110000010100101101010010010011100110001110101100;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b11000110110111000001101111111010110110001111000010111001011101111010110111100010111101010011010011011001001111100100101110111110001111011010110100011001100010011001001100110010011111000110011111011100010100011001100100010111101101000101000111011100110011110000101111010010110100101000101101100100110111011110100111011011111110001100111111011001101110101000101001111110011010011111101001000011100101111100001010000000101101101011100010001000010101001111110001110000111101101110101000000011000000000011100110001011110001011011011100011010111111;
    #1;
    if (!detection)
      failures = failures+1;

    received <= 542'b00111000100101101110100001100000000011110010100000001011100010101001000100001010010011110001101000101001010001101111110101011010000000010001101110111010100010011010111101001110101010001100111111111101111111111000110010001101110110110101110101110000110001000111110101000011001101001001000111000110001000100111001111100011001111110100001111001100001100000010110000011111101100111110010000100011011111101010010101110100001010101110011110001111011010011110101111110101000010101011101010100001100010101001011010010001000100011101011011110001001110;
    #1;
    if (!detection)
      failures = failures+1;

    $display("\n==============================");
    if (!failures)
      $display("\nAll decoding tests passed\n");
    else
      $display("Failed %d decoding test(s)", failures);
    $display("==============================\n");
  end
endmodule
