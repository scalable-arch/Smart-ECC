module bch_encoder(message, codeword);
  input   [511:0] message;
  output  [543:0] codeword;
  wire    [541:0] _codeword;

  assign codeword = {2'b00, 
                    _codeword[29:24], _codeword[541:414], 
                    _codeword[23:16], _codeword[413:286], 
                    _codeword[15:8],  _codeword[285:158], 
                    _codeword[7:0],   _codeword[157:30] };

  assign _codeword[0] = message[0] ^ message[2] ^ message[4] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[10] ^ message[12] ^ message[13] ^ message[14] ^ message[17] ^ message[23] ^ message[24] ^ message[25] ^ message[27] ^ message[28] ^ message[29] ^ message[33] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[42] ^ message[44] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[52] ^ message[54] ^ message[55] ^ message[58] ^ message[60] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[69] ^ message[70] ^ message[73] ^ message[77] ^ message[79] ^ message[81] ^ message[84] ^ message[86] ^ message[88] ^ message[90] ^ message[92] ^ message[93] ^ message[94] ^ message[95] ^ message[97] ^ message[99] ^ message[100] ^ message[101] ^ message[104] ^ message[108] ^ message[109] ^ message[110] ^ message[112] ^ message[114] ^ message[116] ^ message[117] ^ message[120] ^ message[127] ^ message[133] ^ message[135] ^ message[136] ^ message[138] ^ message[139] ^ message[141] ^ message[142] ^ message[146] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[158] ^ message[159] ^ message[161] ^ message[163] ^ message[164] ^ message[166] ^ message[169] ^ message[171] ^ message[173] ^ message[174] ^ message[176] ^ message[177] ^ message[178] ^ message[181] ^ message[183] ^ message[185] ^ message[187] ^ message[189] ^ message[190] ^ message[191] ^ message[194] ^ message[195] ^ message[196] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[214] ^ message[222] ^ message[226] ^ message[228] ^ message[229] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[242] ^ message[244] ^ message[246] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[257] ^ message[258] ^ message[260] ^ message[264] ^ message[265] ^ message[269] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[280] ^ message[282] ^ message[283] ^ message[284] ^ message[294] ^ message[296] ^ message[298] ^ message[300] ^ message[302] ^ message[305] ^ message[309] ^ message[310] ^ message[313] ^ message[315] ^ message[316] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[327] ^ message[329] ^ message[332] ^ message[333] ^ message[334] ^ message[341] ^ message[342] ^ message[343] ^ message[348] ^ message[350] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[360] ^ message[361] ^ message[362] ^ message[363] ^ message[366] ^ message[368] ^ message[369] ^ message[377] ^ message[379] ^ message[380] ^ message[381] ^ message[384] ^ message[385] ^ message[386] ^ message[388] ^ message[389] ^ message[391] ^ message[392] ^ message[393] ^ message[396] ^ message[398] ^ message[400] ^ message[406] ^ message[408] ^ message[409] ^ message[410] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[419] ^ message[420] ^ message[424] ^ message[426] ^ message[429] ^ message[431] ^ message[432] ^ message[433] ^ message[438] ^ message[440] ^ message[442] ^ message[444] ^ message[450] ^ message[451] ^ message[452] ^ message[453] ^ message[455] ^ message[456] ^ message[457] ^ message[459] ^ message[460] ^ message[461] ^ message[472] ^ message[474] ^ message[475] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[485] ^ message[487] ^ message[490] ^ message[492] ^ message[494] ^ message[495] ^ message[496] ^ message[501] ^ message[502] ^ message[503] ^ message[506] ^ message[509];
  assign _codeword[1] = message[0] ^ message[1] ^ message[2] ^ message[3] ^ message[4] ^ message[5] ^ message[6] ^ message[11] ^ message[12] ^ message[15] ^ message[17] ^ message[18] ^ message[23] ^ message[26] ^ message[27] ^ message[30] ^ message[33] ^ message[34] ^ message[35] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[56] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[66] ^ message[69] ^ message[71] ^ message[73] ^ message[74] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[102] ^ message[104] ^ message[105] ^ message[108] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[118] ^ message[120] ^ message[121] ^ message[127] ^ message[128] ^ message[133] ^ message[134] ^ message[135] ^ message[137] ^ message[138] ^ message[140] ^ message[141] ^ message[143] ^ message[146] ^ message[147] ^ message[148] ^ message[153] ^ message[158] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[165] ^ message[166] ^ message[167] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[175] ^ message[176] ^ message[179] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[192] ^ message[194] ^ message[197] ^ message[200] ^ message[206] ^ message[214] ^ message[215] ^ message[222] ^ message[223] ^ message[226] ^ message[227] ^ message[228] ^ message[230] ^ message[231] ^ message[235] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[251] ^ message[255] ^ message[257] ^ message[259] ^ message[260] ^ message[261] ^ message[264] ^ message[266] ^ message[269] ^ message[270] ^ message[272] ^ message[276] ^ message[280] ^ message[281] ^ message[282] ^ message[285] ^ message[294] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[305] ^ message[306] ^ message[309] ^ message[311] ^ message[313] ^ message[314] ^ message[315] ^ message[317] ^ message[320] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[332] ^ message[335] ^ message[341] ^ message[344] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[355] ^ message[359] ^ message[360] ^ message[364] ^ message[366] ^ message[367] ^ message[368] ^ message[370] ^ message[377] ^ message[378] ^ message[379] ^ message[382] ^ message[384] ^ message[387] ^ message[388] ^ message[390] ^ message[391] ^ message[394] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[406] ^ message[407] ^ message[408] ^ message[411] ^ message[412] ^ message[416] ^ message[419] ^ message[421] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[429] ^ message[430] ^ message[431] ^ message[434] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[450] ^ message[454] ^ message[455] ^ message[458] ^ message[459] ^ message[462] ^ message[472] ^ message[473] ^ message[474] ^ message[476] ^ message[478] ^ message[482] ^ message[485] ^ message[486] ^ message[487] ^ message[488] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[497] ^ message[501] ^ message[504] ^ message[506] ^ message[507] ^ message[509] ^ message[510];
  assign _codeword[2] = message[1] ^ message[2] ^ message[3] ^ message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[12] ^ message[13] ^ message[16] ^ message[18] ^ message[19] ^ message[24] ^ message[27] ^ message[28] ^ message[31] ^ message[34] ^ message[35] ^ message[36] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[57] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[67] ^ message[70] ^ message[72] ^ message[74] ^ message[75] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[103] ^ message[105] ^ message[106] ^ message[109] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[119] ^ message[121] ^ message[122] ^ message[128] ^ message[129] ^ message[134] ^ message[135] ^ message[136] ^ message[138] ^ message[139] ^ message[141] ^ message[142] ^ message[144] ^ message[147] ^ message[148] ^ message[149] ^ message[154] ^ message[159] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[166] ^ message[167] ^ message[168] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[176] ^ message[177] ^ message[180] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[193] ^ message[195] ^ message[198] ^ message[201] ^ message[207] ^ message[215] ^ message[216] ^ message[223] ^ message[224] ^ message[227] ^ message[228] ^ message[229] ^ message[231] ^ message[232] ^ message[236] ^ message[243] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[248] ^ message[252] ^ message[256] ^ message[258] ^ message[260] ^ message[261] ^ message[262] ^ message[265] ^ message[267] ^ message[270] ^ message[271] ^ message[273] ^ message[277] ^ message[281] ^ message[282] ^ message[283] ^ message[286] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[306] ^ message[307] ^ message[310] ^ message[312] ^ message[314] ^ message[315] ^ message[316] ^ message[318] ^ message[321] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[333] ^ message[336] ^ message[342] ^ message[345] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[356] ^ message[360] ^ message[361] ^ message[365] ^ message[367] ^ message[368] ^ message[369] ^ message[371] ^ message[378] ^ message[379] ^ message[380] ^ message[383] ^ message[385] ^ message[388] ^ message[389] ^ message[391] ^ message[392] ^ message[395] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[407] ^ message[408] ^ message[409] ^ message[412] ^ message[413] ^ message[417] ^ message[420] ^ message[422] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[430] ^ message[431] ^ message[432] ^ message[435] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[451] ^ message[455] ^ message[456] ^ message[459] ^ message[460] ^ message[463] ^ message[473] ^ message[474] ^ message[475] ^ message[477] ^ message[479] ^ message[483] ^ message[486] ^ message[487] ^ message[488] ^ message[489] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[498] ^ message[502] ^ message[505] ^ message[507] ^ message[508] ^ message[510] ^ message[511];
  assign _codeword[3] = message[2] ^ message[3] ^ message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[13] ^ message[14] ^ message[17] ^ message[19] ^ message[20] ^ message[25] ^ message[28] ^ message[29] ^ message[32] ^ message[35] ^ message[36] ^ message[37] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[53] ^ message[54] ^ message[55] ^ message[56] ^ message[58] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[68] ^ message[71] ^ message[73] ^ message[75] ^ message[76] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[84] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[104] ^ message[106] ^ message[107] ^ message[110] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[120] ^ message[122] ^ message[123] ^ message[129] ^ message[130] ^ message[135] ^ message[136] ^ message[137] ^ message[139] ^ message[140] ^ message[142] ^ message[143] ^ message[145] ^ message[148] ^ message[149] ^ message[150] ^ message[155] ^ message[160] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[167] ^ message[168] ^ message[169] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[177] ^ message[178] ^ message[181] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[194] ^ message[196] ^ message[199] ^ message[202] ^ message[208] ^ message[216] ^ message[217] ^ message[224] ^ message[225] ^ message[228] ^ message[229] ^ message[230] ^ message[232] ^ message[233] ^ message[237] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[253] ^ message[257] ^ message[259] ^ message[261] ^ message[262] ^ message[263] ^ message[266] ^ message[268] ^ message[271] ^ message[272] ^ message[274] ^ message[278] ^ message[282] ^ message[283] ^ message[284] ^ message[287] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[307] ^ message[308] ^ message[311] ^ message[313] ^ message[315] ^ message[316] ^ message[317] ^ message[319] ^ message[322] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[334] ^ message[337] ^ message[343] ^ message[346] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[357] ^ message[361] ^ message[362] ^ message[366] ^ message[368] ^ message[369] ^ message[370] ^ message[372] ^ message[379] ^ message[380] ^ message[381] ^ message[384] ^ message[386] ^ message[389] ^ message[390] ^ message[392] ^ message[393] ^ message[396] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[408] ^ message[409] ^ message[410] ^ message[413] ^ message[414] ^ message[418] ^ message[421] ^ message[423] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[431] ^ message[432] ^ message[433] ^ message[436] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[452] ^ message[456] ^ message[457] ^ message[460] ^ message[461] ^ message[464] ^ message[474] ^ message[475] ^ message[476] ^ message[478] ^ message[480] ^ message[484] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[499] ^ message[503] ^ message[506] ^ message[508] ^ message[509] ^ message[511];
  assign _codeword[4] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[10] ^ message[12] ^ message[13] ^ message[15] ^ message[17] ^ message[18] ^ message[20] ^ message[21] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[30] ^ message[35] ^ message[39] ^ message[40] ^ message[42] ^ message[45] ^ message[50] ^ message[52] ^ message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[70] ^ message[72] ^ message[73] ^ message[74] ^ message[76] ^ message[79] ^ message[80] ^ message[82] ^ message[83] ^ message[85] ^ message[86] ^ message[87] ^ message[89] ^ message[91] ^ message[97] ^ message[102] ^ message[104] ^ message[105] ^ message[107] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[115] ^ message[118] ^ message[119] ^ message[120] ^ message[121] ^ message[123] ^ message[124] ^ message[127] ^ message[130] ^ message[131] ^ message[133] ^ message[135] ^ message[137] ^ message[139] ^ message[140] ^ message[142] ^ message[143] ^ message[144] ^ message[148] ^ message[152] ^ message[156] ^ message[158] ^ message[159] ^ message[165] ^ message[168] ^ message[170] ^ message[171] ^ message[172] ^ message[175] ^ message[177] ^ message[179] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[186] ^ message[188] ^ message[192] ^ message[194] ^ message[196] ^ message[197] ^ message[201] ^ message[202] ^ message[204] ^ message[205] ^ message[209] ^ message[214] ^ message[217] ^ message[218] ^ message[222] ^ message[225] ^ message[228] ^ message[230] ^ message[232] ^ message[238] ^ message[242] ^ message[244] ^ message[245] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[257] ^ message[262] ^ message[263] ^ message[265] ^ message[267] ^ message[274] ^ message[279] ^ message[280] ^ message[282] ^ message[285] ^ message[288] ^ message[294] ^ message[296] ^ message[297] ^ message[299] ^ message[301] ^ message[303] ^ message[304] ^ message[306] ^ message[308] ^ message[310] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[317] ^ message[318] ^ message[321] ^ message[322] ^ message[324] ^ message[325] ^ message[327] ^ message[330] ^ message[331] ^ message[334] ^ message[335] ^ message[338] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[347] ^ message[348] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[360] ^ message[361] ^ message[366] ^ message[367] ^ message[368] ^ message[370] ^ message[371] ^ message[373] ^ message[377] ^ message[379] ^ message[382] ^ message[384] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[392] ^ message[394] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[406] ^ message[408] ^ message[411] ^ message[412] ^ message[413] ^ message[420] ^ message[422] ^ message[426] ^ message[427] ^ message[428] ^ message[430] ^ message[431] ^ message[434] ^ message[437] ^ message[438] ^ message[440] ^ message[441] ^ message[443] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[450] ^ message[451] ^ message[452] ^ message[455] ^ message[456] ^ message[458] ^ message[459] ^ message[460] ^ message[462] ^ message[465] ^ message[472] ^ message[474] ^ message[476] ^ message[477] ^ message[478] ^ message[480] ^ message[487] ^ message[488] ^ message[489] ^ message[491] ^ message[492] ^ message[493] ^ message[497] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[506] ^ message[507] ^ message[510];
  assign _codeword[5] = message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[11] ^ message[13] ^ message[14] ^ message[16] ^ message[18] ^ message[19] ^ message[21] ^ message[22] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[31] ^ message[36] ^ message[40] ^ message[41] ^ message[43] ^ message[46] ^ message[51] ^ message[53] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[71] ^ message[73] ^ message[74] ^ message[75] ^ message[77] ^ message[80] ^ message[81] ^ message[83] ^ message[84] ^ message[86] ^ message[87] ^ message[88] ^ message[90] ^ message[92] ^ message[98] ^ message[103] ^ message[105] ^ message[106] ^ message[108] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[116] ^ message[119] ^ message[120] ^ message[121] ^ message[122] ^ message[124] ^ message[125] ^ message[128] ^ message[131] ^ message[132] ^ message[134] ^ message[136] ^ message[138] ^ message[140] ^ message[141] ^ message[143] ^ message[144] ^ message[145] ^ message[149] ^ message[153] ^ message[157] ^ message[159] ^ message[160] ^ message[166] ^ message[169] ^ message[171] ^ message[172] ^ message[173] ^ message[176] ^ message[178] ^ message[180] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[187] ^ message[189] ^ message[193] ^ message[195] ^ message[197] ^ message[198] ^ message[202] ^ message[203] ^ message[205] ^ message[206] ^ message[210] ^ message[215] ^ message[218] ^ message[219] ^ message[223] ^ message[226] ^ message[229] ^ message[231] ^ message[233] ^ message[239] ^ message[243] ^ message[245] ^ message[246] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[258] ^ message[263] ^ message[264] ^ message[266] ^ message[268] ^ message[275] ^ message[280] ^ message[281] ^ message[283] ^ message[286] ^ message[289] ^ message[295] ^ message[297] ^ message[298] ^ message[300] ^ message[302] ^ message[304] ^ message[305] ^ message[307] ^ message[309] ^ message[311] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[318] ^ message[319] ^ message[322] ^ message[323] ^ message[325] ^ message[326] ^ message[328] ^ message[331] ^ message[332] ^ message[335] ^ message[336] ^ message[339] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[348] ^ message[349] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[361] ^ message[362] ^ message[367] ^ message[368] ^ message[369] ^ message[371] ^ message[372] ^ message[374] ^ message[378] ^ message[380] ^ message[383] ^ message[385] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[393] ^ message[395] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[407] ^ message[409] ^ message[412] ^ message[413] ^ message[414] ^ message[421] ^ message[423] ^ message[427] ^ message[428] ^ message[429] ^ message[431] ^ message[432] ^ message[435] ^ message[438] ^ message[439] ^ message[441] ^ message[442] ^ message[444] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[451] ^ message[452] ^ message[453] ^ message[456] ^ message[457] ^ message[459] ^ message[460] ^ message[461] ^ message[463] ^ message[466] ^ message[473] ^ message[475] ^ message[477] ^ message[478] ^ message[479] ^ message[481] ^ message[488] ^ message[489] ^ message[490] ^ message[492] ^ message[493] ^ message[494] ^ message[498] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[507] ^ message[508] ^ message[511];
  assign _codeword[6] = message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[12] ^ message[14] ^ message[15] ^ message[17] ^ message[19] ^ message[20] ^ message[22] ^ message[23] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[32] ^ message[37] ^ message[41] ^ message[42] ^ message[44] ^ message[47] ^ message[52] ^ message[54] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[72] ^ message[74] ^ message[75] ^ message[76] ^ message[78] ^ message[81] ^ message[82] ^ message[84] ^ message[85] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[93] ^ message[99] ^ message[104] ^ message[106] ^ message[107] ^ message[109] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[117] ^ message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[125] ^ message[126] ^ message[129] ^ message[132] ^ message[133] ^ message[135] ^ message[137] ^ message[139] ^ message[141] ^ message[142] ^ message[144] ^ message[145] ^ message[146] ^ message[150] ^ message[154] ^ message[158] ^ message[160] ^ message[161] ^ message[167] ^ message[170] ^ message[172] ^ message[173] ^ message[174] ^ message[177] ^ message[179] ^ message[181] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[188] ^ message[190] ^ message[194] ^ message[196] ^ message[198] ^ message[199] ^ message[203] ^ message[204] ^ message[206] ^ message[207] ^ message[211] ^ message[216] ^ message[219] ^ message[220] ^ message[224] ^ message[227] ^ message[230] ^ message[232] ^ message[234] ^ message[240] ^ message[244] ^ message[246] ^ message[247] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[259] ^ message[264] ^ message[265] ^ message[267] ^ message[269] ^ message[276] ^ message[281] ^ message[282] ^ message[284] ^ message[287] ^ message[290] ^ message[296] ^ message[298] ^ message[299] ^ message[301] ^ message[303] ^ message[305] ^ message[306] ^ message[308] ^ message[310] ^ message[312] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[319] ^ message[320] ^ message[323] ^ message[324] ^ message[326] ^ message[327] ^ message[329] ^ message[332] ^ message[333] ^ message[336] ^ message[337] ^ message[340] ^ message[343] ^ message[344] ^ message[345] ^ message[346] ^ message[349] ^ message[350] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[362] ^ message[363] ^ message[368] ^ message[369] ^ message[370] ^ message[372] ^ message[373] ^ message[375] ^ message[379] ^ message[381] ^ message[384] ^ message[386] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[394] ^ message[396] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[408] ^ message[410] ^ message[413] ^ message[414] ^ message[415] ^ message[422] ^ message[424] ^ message[428] ^ message[429] ^ message[430] ^ message[432] ^ message[433] ^ message[436] ^ message[439] ^ message[440] ^ message[442] ^ message[443] ^ message[445] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[452] ^ message[453] ^ message[454] ^ message[457] ^ message[458] ^ message[460] ^ message[461] ^ message[462] ^ message[464] ^ message[467] ^ message[474] ^ message[476] ^ message[478] ^ message[479] ^ message[480] ^ message[482] ^ message[489] ^ message[490] ^ message[491] ^ message[493] ^ message[494] ^ message[495] ^ message[499] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[508] ^ message[509];
  assign _codeword[7] = message[3] ^ message[5] ^ message[6] ^ message[8] ^ message[13] ^ message[15] ^ message[16] ^ message[18] ^ message[20] ^ message[21] ^ message[23] ^ message[24] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[33] ^ message[38] ^ message[42] ^ message[43] ^ message[45] ^ message[48] ^ message[53] ^ message[55] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[73] ^ message[75] ^ message[76] ^ message[77] ^ message[79] ^ message[82] ^ message[83] ^ message[85] ^ message[86] ^ message[88] ^ message[89] ^ message[90] ^ message[92] ^ message[94] ^ message[100] ^ message[105] ^ message[107] ^ message[108] ^ message[110] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[118] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[126] ^ message[127] ^ message[130] ^ message[133] ^ message[134] ^ message[136] ^ message[138] ^ message[140] ^ message[142] ^ message[143] ^ message[145] ^ message[146] ^ message[147] ^ message[151] ^ message[155] ^ message[159] ^ message[161] ^ message[162] ^ message[168] ^ message[171] ^ message[173] ^ message[174] ^ message[175] ^ message[178] ^ message[180] ^ message[182] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[189] ^ message[191] ^ message[195] ^ message[197] ^ message[199] ^ message[200] ^ message[204] ^ message[205] ^ message[207] ^ message[208] ^ message[212] ^ message[217] ^ message[220] ^ message[221] ^ message[225] ^ message[228] ^ message[231] ^ message[233] ^ message[235] ^ message[241] ^ message[245] ^ message[247] ^ message[248] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[256] ^ message[260] ^ message[265] ^ message[266] ^ message[268] ^ message[270] ^ message[277] ^ message[282] ^ message[283] ^ message[285] ^ message[288] ^ message[291] ^ message[297] ^ message[299] ^ message[300] ^ message[302] ^ message[304] ^ message[306] ^ message[307] ^ message[309] ^ message[311] ^ message[313] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[320] ^ message[321] ^ message[324] ^ message[325] ^ message[327] ^ message[328] ^ message[330] ^ message[333] ^ message[334] ^ message[337] ^ message[338] ^ message[341] ^ message[344] ^ message[345] ^ message[346] ^ message[347] ^ message[350] ^ message[351] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[363] ^ message[364] ^ message[369] ^ message[370] ^ message[371] ^ message[373] ^ message[374] ^ message[376] ^ message[380] ^ message[382] ^ message[385] ^ message[387] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[395] ^ message[397] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[409] ^ message[411] ^ message[414] ^ message[415] ^ message[416] ^ message[423] ^ message[425] ^ message[429] ^ message[430] ^ message[431] ^ message[433] ^ message[434] ^ message[437] ^ message[440] ^ message[441] ^ message[443] ^ message[444] ^ message[446] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[453] ^ message[454] ^ message[455] ^ message[458] ^ message[459] ^ message[461] ^ message[462] ^ message[463] ^ message[465] ^ message[468] ^ message[475] ^ message[477] ^ message[479] ^ message[480] ^ message[481] ^ message[483] ^ message[490] ^ message[491] ^ message[492] ^ message[494] ^ message[495] ^ message[496] ^ message[500] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[507] ^ message[509] ^ message[510];
  assign _codeword[8] = message[0] ^ message[2] ^ message[8] ^ message[10] ^ message[12] ^ message[13] ^ message[16] ^ message[19] ^ message[21] ^ message[22] ^ message[23] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[40] ^ message[42] ^ message[43] ^ message[47] ^ message[48] ^ message[50] ^ message[52] ^ message[55] ^ message[56] ^ message[58] ^ message[61] ^ message[69] ^ message[70] ^ message[73] ^ message[74] ^ message[76] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[83] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[92] ^ message[94] ^ message[97] ^ message[99] ^ message[100] ^ message[104] ^ message[106] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[115] ^ message[117] ^ message[119] ^ message[120] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[128] ^ message[131] ^ message[133] ^ message[134] ^ message[136] ^ message[137] ^ message[138] ^ message[142] ^ message[143] ^ message[144] ^ message[147] ^ message[149] ^ message[150] ^ message[151] ^ message[156] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[164] ^ message[166] ^ message[171] ^ message[172] ^ message[173] ^ message[175] ^ message[177] ^ message[178] ^ message[179] ^ message[186] ^ message[188] ^ message[189] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[198] ^ message[202] ^ message[203] ^ message[204] ^ message[206] ^ message[208] ^ message[209] ^ message[213] ^ message[214] ^ message[218] ^ message[221] ^ message[228] ^ message[231] ^ message[233] ^ message[236] ^ message[244] ^ message[248] ^ message[249] ^ message[255] ^ message[256] ^ message[258] ^ message[260] ^ message[261] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[278] ^ message[280] ^ message[282] ^ message[286] ^ message[289] ^ message[292] ^ message[294] ^ message[296] ^ message[301] ^ message[302] ^ message[303] ^ message[307] ^ message[308] ^ message[309] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[323] ^ message[324] ^ message[326] ^ message[327] ^ message[328] ^ message[331] ^ message[332] ^ message[333] ^ message[335] ^ message[338] ^ message[339] ^ message[341] ^ message[343] ^ message[345] ^ message[346] ^ message[347] ^ message[350] ^ message[351] ^ message[352] ^ message[354] ^ message[359] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[368] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[374] ^ message[375] ^ message[379] ^ message[380] ^ message[383] ^ message[384] ^ message[385] ^ message[389] ^ message[390] ^ message[394] ^ message[401] ^ message[402] ^ message[403] ^ message[405] ^ message[407] ^ message[409] ^ message[413] ^ message[414] ^ message[416] ^ message[417] ^ message[419] ^ message[420] ^ message[429] ^ message[430] ^ message[433] ^ message[434] ^ message[435] ^ message[440] ^ message[441] ^ message[445] ^ message[447] ^ message[449] ^ message[453] ^ message[454] ^ message[457] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[466] ^ message[469] ^ message[472] ^ message[474] ^ message[475] ^ message[476] ^ message[479] ^ message[482] ^ message[484] ^ message[485] ^ message[487] ^ message[490] ^ message[491] ^ message[493] ^ message[494] ^ message[497] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511];
  assign _codeword[9] = message[1] ^ message[3] ^ message[9] ^ message[11] ^ message[13] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[23] ^ message[24] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[41] ^ message[43] ^ message[44] ^ message[48] ^ message[49] ^ message[51] ^ message[53] ^ message[56] ^ message[57] ^ message[59] ^ message[62] ^ message[70] ^ message[71] ^ message[74] ^ message[75] ^ message[77] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[84] ^ message[88] ^ message[89] ^ message[90] ^ message[92] ^ message[93] ^ message[95] ^ message[98] ^ message[100] ^ message[101] ^ message[105] ^ message[107] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[116] ^ message[118] ^ message[120] ^ message[121] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[129] ^ message[132] ^ message[134] ^ message[135] ^ message[137] ^ message[138] ^ message[139] ^ message[143] ^ message[144] ^ message[145] ^ message[148] ^ message[150] ^ message[151] ^ message[152] ^ message[157] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[165] ^ message[167] ^ message[172] ^ message[173] ^ message[174] ^ message[176] ^ message[178] ^ message[179] ^ message[180] ^ message[187] ^ message[189] ^ message[190] ^ message[192] ^ message[193] ^ message[195] ^ message[196] ^ message[199] ^ message[203] ^ message[204] ^ message[205] ^ message[207] ^ message[209] ^ message[210] ^ message[214] ^ message[215] ^ message[219] ^ message[222] ^ message[229] ^ message[232] ^ message[234] ^ message[237] ^ message[245] ^ message[249] ^ message[250] ^ message[256] ^ message[257] ^ message[259] ^ message[261] ^ message[262] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[279] ^ message[281] ^ message[283] ^ message[287] ^ message[290] ^ message[293] ^ message[295] ^ message[297] ^ message[302] ^ message[303] ^ message[304] ^ message[308] ^ message[309] ^ message[310] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[324] ^ message[325] ^ message[327] ^ message[328] ^ message[329] ^ message[332] ^ message[333] ^ message[334] ^ message[336] ^ message[339] ^ message[340] ^ message[342] ^ message[344] ^ message[346] ^ message[347] ^ message[348] ^ message[351] ^ message[352] ^ message[353] ^ message[355] ^ message[360] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[375] ^ message[376] ^ message[380] ^ message[381] ^ message[384] ^ message[385] ^ message[386] ^ message[390] ^ message[391] ^ message[395] ^ message[402] ^ message[403] ^ message[404] ^ message[406] ^ message[408] ^ message[410] ^ message[414] ^ message[415] ^ message[417] ^ message[418] ^ message[420] ^ message[421] ^ message[430] ^ message[431] ^ message[434] ^ message[435] ^ message[436] ^ message[441] ^ message[442] ^ message[446] ^ message[448] ^ message[450] ^ message[454] ^ message[455] ^ message[458] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[467] ^ message[470] ^ message[473] ^ message[475] ^ message[476] ^ message[477] ^ message[480] ^ message[483] ^ message[485] ^ message[486] ^ message[488] ^ message[491] ^ message[492] ^ message[494] ^ message[495] ^ message[498] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[508] ^ message[509] ^ message[510] ^ message[511];
  assign _codeword[10] = message[2] ^ message[4] ^ message[10] ^ message[12] ^ message[14] ^ message[15] ^ message[18] ^ message[21] ^ message[23] ^ message[24] ^ message[25] ^ message[32] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[42] ^ message[44] ^ message[45] ^ message[49] ^ message[50] ^ message[52] ^ message[54] ^ message[57] ^ message[58] ^ message[60] ^ message[63] ^ message[71] ^ message[72] ^ message[75] ^ message[76] ^ message[78] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[85] ^ message[89] ^ message[90] ^ message[91] ^ message[93] ^ message[94] ^ message[96] ^ message[99] ^ message[101] ^ message[102] ^ message[106] ^ message[108] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[117] ^ message[119] ^ message[121] ^ message[122] ^ message[124] ^ message[125] ^ message[126] ^ message[127] ^ message[130] ^ message[133] ^ message[135] ^ message[136] ^ message[138] ^ message[139] ^ message[140] ^ message[144] ^ message[145] ^ message[146] ^ message[149] ^ message[151] ^ message[152] ^ message[153] ^ message[158] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[166] ^ message[168] ^ message[173] ^ message[174] ^ message[175] ^ message[177] ^ message[179] ^ message[180] ^ message[181] ^ message[188] ^ message[190] ^ message[191] ^ message[193] ^ message[194] ^ message[196] ^ message[197] ^ message[200] ^ message[204] ^ message[205] ^ message[206] ^ message[208] ^ message[210] ^ message[211] ^ message[215] ^ message[216] ^ message[220] ^ message[223] ^ message[230] ^ message[233] ^ message[235] ^ message[238] ^ message[246] ^ message[250] ^ message[251] ^ message[257] ^ message[258] ^ message[260] ^ message[262] ^ message[263] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[280] ^ message[282] ^ message[284] ^ message[288] ^ message[291] ^ message[294] ^ message[296] ^ message[298] ^ message[303] ^ message[304] ^ message[305] ^ message[309] ^ message[310] ^ message[311] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[325] ^ message[326] ^ message[328] ^ message[329] ^ message[330] ^ message[333] ^ message[334] ^ message[335] ^ message[337] ^ message[340] ^ message[341] ^ message[343] ^ message[345] ^ message[347] ^ message[348] ^ message[349] ^ message[352] ^ message[353] ^ message[354] ^ message[356] ^ message[361] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[376] ^ message[377] ^ message[381] ^ message[382] ^ message[385] ^ message[386] ^ message[387] ^ message[391] ^ message[392] ^ message[396] ^ message[403] ^ message[404] ^ message[405] ^ message[407] ^ message[409] ^ message[411] ^ message[415] ^ message[416] ^ message[418] ^ message[419] ^ message[421] ^ message[422] ^ message[431] ^ message[432] ^ message[435] ^ message[436] ^ message[437] ^ message[442] ^ message[443] ^ message[447] ^ message[449] ^ message[451] ^ message[455] ^ message[456] ^ message[459] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[468] ^ message[471] ^ message[474] ^ message[476] ^ message[477] ^ message[478] ^ message[481] ^ message[484] ^ message[486] ^ message[487] ^ message[489] ^ message[492] ^ message[493] ^ message[495] ^ message[496] ^ message[499] ^ message[504] ^ message[505] ^ message[506] ^ message[507] ^ message[509] ^ message[510] ^ message[511];
  assign _codeword[11] = message[3] ^ message[5] ^ message[11] ^ message[13] ^ message[15] ^ message[16] ^ message[19] ^ message[22] ^ message[24] ^ message[25] ^ message[26] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[43] ^ message[45] ^ message[46] ^ message[50] ^ message[51] ^ message[53] ^ message[55] ^ message[58] ^ message[59] ^ message[61] ^ message[64] ^ message[72] ^ message[73] ^ message[76] ^ message[77] ^ message[79] ^ message[81] ^ message[82] ^ message[83] ^ message[84] ^ message[86] ^ message[90] ^ message[91] ^ message[92] ^ message[94] ^ message[95] ^ message[97] ^ message[100] ^ message[102] ^ message[103] ^ message[107] ^ message[109] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[118] ^ message[120] ^ message[122] ^ message[123] ^ message[125] ^ message[126] ^ message[127] ^ message[128] ^ message[131] ^ message[134] ^ message[136] ^ message[137] ^ message[139] ^ message[140] ^ message[141] ^ message[145] ^ message[146] ^ message[147] ^ message[150] ^ message[152] ^ message[153] ^ message[154] ^ message[159] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[167] ^ message[169] ^ message[174] ^ message[175] ^ message[176] ^ message[178] ^ message[180] ^ message[181] ^ message[182] ^ message[189] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[197] ^ message[198] ^ message[201] ^ message[205] ^ message[206] ^ message[207] ^ message[209] ^ message[211] ^ message[212] ^ message[216] ^ message[217] ^ message[221] ^ message[224] ^ message[231] ^ message[234] ^ message[236] ^ message[239] ^ message[247] ^ message[251] ^ message[252] ^ message[258] ^ message[259] ^ message[261] ^ message[263] ^ message[264] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[278] ^ message[281] ^ message[283] ^ message[285] ^ message[289] ^ message[292] ^ message[295] ^ message[297] ^ message[299] ^ message[304] ^ message[305] ^ message[306] ^ message[310] ^ message[311] ^ message[312] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[326] ^ message[327] ^ message[329] ^ message[330] ^ message[331] ^ message[334] ^ message[335] ^ message[336] ^ message[338] ^ message[341] ^ message[342] ^ message[344] ^ message[346] ^ message[348] ^ message[349] ^ message[350] ^ message[353] ^ message[354] ^ message[355] ^ message[357] ^ message[362] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[377] ^ message[378] ^ message[382] ^ message[383] ^ message[386] ^ message[387] ^ message[388] ^ message[392] ^ message[393] ^ message[397] ^ message[404] ^ message[405] ^ message[406] ^ message[408] ^ message[410] ^ message[412] ^ message[416] ^ message[417] ^ message[419] ^ message[420] ^ message[422] ^ message[423] ^ message[432] ^ message[433] ^ message[436] ^ message[437] ^ message[438] ^ message[443] ^ message[444] ^ message[448] ^ message[450] ^ message[452] ^ message[456] ^ message[457] ^ message[460] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[469] ^ message[472] ^ message[475] ^ message[477] ^ message[478] ^ message[479] ^ message[482] ^ message[485] ^ message[487] ^ message[488] ^ message[490] ^ message[493] ^ message[494] ^ message[496] ^ message[497] ^ message[500] ^ message[505] ^ message[506] ^ message[507] ^ message[508] ^ message[510] ^ message[511];
  assign _codeword[12] = message[0] ^ message[2] ^ message[7] ^ message[8] ^ message[9] ^ message[10] ^ message[13] ^ message[16] ^ message[20] ^ message[24] ^ message[26] ^ message[28] ^ message[29] ^ message[33] ^ message[34] ^ message[41] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[55] ^ message[56] ^ message[58] ^ message[59] ^ message[63] ^ message[64] ^ message[69] ^ message[70] ^ message[74] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[90] ^ message[91] ^ message[94] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[103] ^ message[109] ^ message[112] ^ message[115] ^ message[119] ^ message[120] ^ message[121] ^ message[123] ^ message[124] ^ message[126] ^ message[128] ^ message[129] ^ message[132] ^ message[133] ^ message[136] ^ message[137] ^ message[139] ^ message[140] ^ message[147] ^ message[149] ^ message[150] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[165] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[173] ^ message[174] ^ message[175] ^ message[178] ^ message[179] ^ message[182] ^ message[185] ^ message[187] ^ message[189] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[210] ^ message[212] ^ message[213] ^ message[214] ^ message[217] ^ message[218] ^ message[225] ^ message[226] ^ message[228] ^ message[229] ^ message[231] ^ message[233] ^ message[234] ^ message[235] ^ message[237] ^ message[240] ^ message[242] ^ message[244] ^ message[246] ^ message[248] ^ message[251] ^ message[254] ^ message[257] ^ message[258] ^ message[259] ^ message[262] ^ message[268] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[283] ^ message[286] ^ message[290] ^ message[293] ^ message[294] ^ message[302] ^ message[306] ^ message[307] ^ message[309] ^ message[310] ^ message[311] ^ message[312] ^ message[315] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[325] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[339] ^ message[341] ^ message[345] ^ message[347] ^ message[348] ^ message[349] ^ message[351] ^ message[354] ^ message[357] ^ message[360] ^ message[361] ^ message[362] ^ message[367] ^ message[370] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[380] ^ message[381] ^ message[383] ^ message[385] ^ message[386] ^ message[387] ^ message[391] ^ message[392] ^ message[394] ^ message[396] ^ message[400] ^ message[405] ^ message[407] ^ message[408] ^ message[410] ^ message[411] ^ message[412] ^ message[414] ^ message[415] ^ message[417] ^ message[418] ^ message[419] ^ message[421] ^ message[423] ^ message[426] ^ message[429] ^ message[431] ^ message[432] ^ message[434] ^ message[437] ^ message[439] ^ message[440] ^ message[442] ^ message[445] ^ message[449] ^ message[450] ^ message[452] ^ message[455] ^ message[456] ^ message[458] ^ message[459] ^ message[460] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[470] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[481] ^ message[483] ^ message[485] ^ message[486] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[496] ^ message[497] ^ message[498] ^ message[502] ^ message[503] ^ message[507] ^ message[508] ^ message[511];
  assign _codeword[13] = message[1] ^ message[3] ^ message[8] ^ message[9] ^ message[10] ^ message[11] ^ message[14] ^ message[17] ^ message[21] ^ message[25] ^ message[27] ^ message[29] ^ message[30] ^ message[34] ^ message[35] ^ message[42] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[56] ^ message[57] ^ message[59] ^ message[60] ^ message[64] ^ message[65] ^ message[70] ^ message[71] ^ message[75] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[84] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[92] ^ message[95] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[104] ^ message[110] ^ message[113] ^ message[116] ^ message[120] ^ message[121] ^ message[122] ^ message[124] ^ message[125] ^ message[127] ^ message[129] ^ message[130] ^ message[133] ^ message[134] ^ message[137] ^ message[138] ^ message[140] ^ message[141] ^ message[148] ^ message[150] ^ message[151] ^ message[153] ^ message[154] ^ message[155] ^ message[156] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[166] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[174] ^ message[175] ^ message[176] ^ message[179] ^ message[180] ^ message[183] ^ message[186] ^ message[188] ^ message[190] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[211] ^ message[213] ^ message[214] ^ message[215] ^ message[218] ^ message[219] ^ message[226] ^ message[227] ^ message[229] ^ message[230] ^ message[232] ^ message[234] ^ message[235] ^ message[236] ^ message[238] ^ message[241] ^ message[243] ^ message[245] ^ message[247] ^ message[249] ^ message[252] ^ message[255] ^ message[258] ^ message[259] ^ message[260] ^ message[263] ^ message[269] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[284] ^ message[287] ^ message[291] ^ message[294] ^ message[295] ^ message[303] ^ message[307] ^ message[308] ^ message[310] ^ message[311] ^ message[312] ^ message[313] ^ message[316] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[326] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[340] ^ message[342] ^ message[346] ^ message[348] ^ message[349] ^ message[350] ^ message[352] ^ message[355] ^ message[358] ^ message[361] ^ message[362] ^ message[363] ^ message[368] ^ message[371] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[381] ^ message[382] ^ message[384] ^ message[386] ^ message[387] ^ message[388] ^ message[392] ^ message[393] ^ message[395] ^ message[397] ^ message[401] ^ message[406] ^ message[408] ^ message[409] ^ message[411] ^ message[412] ^ message[413] ^ message[415] ^ message[416] ^ message[418] ^ message[419] ^ message[420] ^ message[422] ^ message[424] ^ message[427] ^ message[430] ^ message[432] ^ message[433] ^ message[435] ^ message[438] ^ message[440] ^ message[441] ^ message[443] ^ message[446] ^ message[450] ^ message[451] ^ message[453] ^ message[456] ^ message[457] ^ message[459] ^ message[460] ^ message[461] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[471] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[482] ^ message[484] ^ message[486] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[497] ^ message[498] ^ message[499] ^ message[503] ^ message[504] ^ message[508] ^ message[509];
  assign _codeword[14] = message[2] ^ message[4] ^ message[9] ^ message[10] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[22] ^ message[26] ^ message[28] ^ message[30] ^ message[31] ^ message[35] ^ message[36] ^ message[43] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[57] ^ message[58] ^ message[60] ^ message[61] ^ message[65] ^ message[66] ^ message[71] ^ message[72] ^ message[76] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[84] ^ message[85] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[92] ^ message[93] ^ message[96] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[105] ^ message[111] ^ message[114] ^ message[117] ^ message[121] ^ message[122] ^ message[123] ^ message[125] ^ message[126] ^ message[128] ^ message[130] ^ message[131] ^ message[134] ^ message[135] ^ message[138] ^ message[139] ^ message[141] ^ message[142] ^ message[149] ^ message[151] ^ message[152] ^ message[154] ^ message[155] ^ message[156] ^ message[157] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[167] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[175] ^ message[176] ^ message[177] ^ message[180] ^ message[181] ^ message[184] ^ message[187] ^ message[189] ^ message[191] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[212] ^ message[214] ^ message[215] ^ message[216] ^ message[219] ^ message[220] ^ message[227] ^ message[228] ^ message[230] ^ message[231] ^ message[233] ^ message[235] ^ message[236] ^ message[237] ^ message[239] ^ message[242] ^ message[244] ^ message[246] ^ message[248] ^ message[250] ^ message[253] ^ message[256] ^ message[259] ^ message[260] ^ message[261] ^ message[264] ^ message[270] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[285] ^ message[288] ^ message[292] ^ message[295] ^ message[296] ^ message[304] ^ message[308] ^ message[309] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[317] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[327] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[341] ^ message[343] ^ message[347] ^ message[349] ^ message[350] ^ message[351] ^ message[353] ^ message[356] ^ message[359] ^ message[362] ^ message[363] ^ message[364] ^ message[369] ^ message[372] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[382] ^ message[383] ^ message[385] ^ message[387] ^ message[388] ^ message[389] ^ message[393] ^ message[394] ^ message[396] ^ message[398] ^ message[402] ^ message[407] ^ message[409] ^ message[410] ^ message[412] ^ message[413] ^ message[414] ^ message[416] ^ message[417] ^ message[419] ^ message[420] ^ message[421] ^ message[423] ^ message[425] ^ message[428] ^ message[431] ^ message[433] ^ message[434] ^ message[436] ^ message[439] ^ message[441] ^ message[442] ^ message[444] ^ message[447] ^ message[451] ^ message[452] ^ message[454] ^ message[457] ^ message[458] ^ message[460] ^ message[461] ^ message[462] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[472] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[483] ^ message[485] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[498] ^ message[499] ^ message[500] ^ message[504] ^ message[505] ^ message[509] ^ message[510];
  assign _codeword[15] = message[3] ^ message[5] ^ message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[16] ^ message[19] ^ message[23] ^ message[27] ^ message[29] ^ message[31] ^ message[32] ^ message[36] ^ message[37] ^ message[44] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[58] ^ message[59] ^ message[61] ^ message[62] ^ message[66] ^ message[67] ^ message[72] ^ message[73] ^ message[77] ^ message[81] ^ message[82] ^ message[83] ^ message[84] ^ message[85] ^ message[86] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[93] ^ message[94] ^ message[97] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[106] ^ message[112] ^ message[115] ^ message[118] ^ message[122] ^ message[123] ^ message[124] ^ message[126] ^ message[127] ^ message[129] ^ message[131] ^ message[132] ^ message[135] ^ message[136] ^ message[139] ^ message[140] ^ message[142] ^ message[143] ^ message[150] ^ message[152] ^ message[153] ^ message[155] ^ message[156] ^ message[157] ^ message[158] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[168] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[176] ^ message[177] ^ message[178] ^ message[181] ^ message[182] ^ message[185] ^ message[188] ^ message[190] ^ message[192] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[213] ^ message[215] ^ message[216] ^ message[217] ^ message[220] ^ message[221] ^ message[228] ^ message[229] ^ message[231] ^ message[232] ^ message[234] ^ message[236] ^ message[237] ^ message[238] ^ message[240] ^ message[243] ^ message[245] ^ message[247] ^ message[249] ^ message[251] ^ message[254] ^ message[257] ^ message[260] ^ message[261] ^ message[262] ^ message[265] ^ message[271] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[283] ^ message[286] ^ message[289] ^ message[293] ^ message[296] ^ message[297] ^ message[305] ^ message[309] ^ message[310] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[318] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[328] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[342] ^ message[344] ^ message[348] ^ message[350] ^ message[351] ^ message[352] ^ message[354] ^ message[357] ^ message[360] ^ message[363] ^ message[364] ^ message[365] ^ message[370] ^ message[373] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[381] ^ message[383] ^ message[384] ^ message[386] ^ message[388] ^ message[389] ^ message[390] ^ message[394] ^ message[395] ^ message[397] ^ message[399] ^ message[403] ^ message[408] ^ message[410] ^ message[411] ^ message[413] ^ message[414] ^ message[415] ^ message[417] ^ message[418] ^ message[420] ^ message[421] ^ message[422] ^ message[424] ^ message[426] ^ message[429] ^ message[432] ^ message[434] ^ message[435] ^ message[437] ^ message[440] ^ message[442] ^ message[443] ^ message[445] ^ message[448] ^ message[452] ^ message[453] ^ message[455] ^ message[458] ^ message[459] ^ message[461] ^ message[462] ^ message[463] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[473] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[484] ^ message[486] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[499] ^ message[500] ^ message[501] ^ message[505] ^ message[506] ^ message[510] ^ message[511];
  assign _codeword[16] = message[0] ^ message[2] ^ message[7] ^ message[8] ^ message[9] ^ message[10] ^ message[11] ^ message[20] ^ message[23] ^ message[25] ^ message[27] ^ message[29] ^ message[30] ^ message[32] ^ message[35] ^ message[36] ^ message[39] ^ message[40] ^ message[42] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[53] ^ message[58] ^ message[59] ^ message[64] ^ message[65] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[74] ^ message[77] ^ message[78] ^ message[79] ^ message[81] ^ message[82] ^ message[83] ^ message[85] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[93] ^ message[97] ^ message[98] ^ message[99] ^ message[102] ^ message[103] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[112] ^ message[113] ^ message[114] ^ message[117] ^ message[119] ^ message[120] ^ message[123] ^ message[124] ^ message[125] ^ message[128] ^ message[130] ^ message[132] ^ message[135] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[142] ^ message[143] ^ message[144] ^ message[146] ^ message[148] ^ message[149] ^ message[150] ^ message[152] ^ message[153] ^ message[154] ^ message[156] ^ message[157] ^ message[161] ^ message[162] ^ message[165] ^ message[171] ^ message[172] ^ message[175] ^ message[176] ^ message[179] ^ message[181] ^ message[182] ^ message[185] ^ message[186] ^ message[187] ^ message[190] ^ message[193] ^ message[194] ^ message[197] ^ message[198] ^ message[200] ^ message[201] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[216] ^ message[217] ^ message[218] ^ message[221] ^ message[226] ^ message[228] ^ message[230] ^ message[231] ^ message[234] ^ message[235] ^ message[237] ^ message[238] ^ message[239] ^ message[241] ^ message[242] ^ message[248] ^ message[250] ^ message[251] ^ message[253] ^ message[254] ^ message[255] ^ message[257] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[269] ^ message[273] ^ message[276] ^ message[277] ^ message[278] ^ message[281] ^ message[287] ^ message[290] ^ message[296] ^ message[297] ^ message[300] ^ message[302] ^ message[305] ^ message[306] ^ message[309] ^ message[311] ^ message[314] ^ message[319] ^ message[320] ^ message[325] ^ message[327] ^ message[335] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[342] ^ message[345] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[356] ^ message[357] ^ message[360] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[368] ^ message[369] ^ message[371] ^ message[374] ^ message[376] ^ message[378] ^ message[382] ^ message[386] ^ message[387] ^ message[388] ^ message[390] ^ message[392] ^ message[393] ^ message[395] ^ message[404] ^ message[406] ^ message[408] ^ message[410] ^ message[411] ^ message[413] ^ message[416] ^ message[418] ^ message[420] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[429] ^ message[430] ^ message[431] ^ message[432] ^ message[435] ^ message[436] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[446] ^ message[449] ^ message[450] ^ message[451] ^ message[452] ^ message[454] ^ message[455] ^ message[457] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[469] ^ message[470] ^ message[471] ^ message[475] ^ message[476] ^ message[477] ^ message[481] ^ message[489] ^ message[491] ^ message[493] ^ message[500] ^ message[503] ^ message[507] ^ message[509] ^ message[511];
  assign _codeword[17] = message[1] ^ message[3] ^ message[8] ^ message[9] ^ message[10] ^ message[11] ^ message[12] ^ message[21] ^ message[24] ^ message[26] ^ message[28] ^ message[30] ^ message[31] ^ message[33] ^ message[36] ^ message[37] ^ message[40] ^ message[41] ^ message[43] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[54] ^ message[59] ^ message[60] ^ message[65] ^ message[66] ^ message[68] ^ message[69] ^ message[70] ^ message[71] ^ message[75] ^ message[78] ^ message[79] ^ message[80] ^ message[82] ^ message[83] ^ message[84] ^ message[86] ^ message[88] ^ message[89] ^ message[90] ^ message[92] ^ message[94] ^ message[98] ^ message[99] ^ message[100] ^ message[103] ^ message[104] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[113] ^ message[114] ^ message[115] ^ message[118] ^ message[120] ^ message[121] ^ message[124] ^ message[125] ^ message[126] ^ message[129] ^ message[131] ^ message[133] ^ message[136] ^ message[138] ^ message[139] ^ message[140] ^ message[141] ^ message[143] ^ message[144] ^ message[145] ^ message[147] ^ message[149] ^ message[150] ^ message[151] ^ message[153] ^ message[154] ^ message[155] ^ message[157] ^ message[158] ^ message[162] ^ message[163] ^ message[166] ^ message[172] ^ message[173] ^ message[176] ^ message[177] ^ message[180] ^ message[182] ^ message[183] ^ message[186] ^ message[187] ^ message[188] ^ message[191] ^ message[194] ^ message[195] ^ message[198] ^ message[199] ^ message[201] ^ message[202] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[217] ^ message[218] ^ message[219] ^ message[222] ^ message[227] ^ message[229] ^ message[231] ^ message[232] ^ message[235] ^ message[236] ^ message[238] ^ message[239] ^ message[240] ^ message[242] ^ message[243] ^ message[249] ^ message[251] ^ message[252] ^ message[254] ^ message[255] ^ message[256] ^ message[258] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[270] ^ message[274] ^ message[277] ^ message[278] ^ message[279] ^ message[282] ^ message[288] ^ message[291] ^ message[297] ^ message[298] ^ message[301] ^ message[303] ^ message[306] ^ message[307] ^ message[310] ^ message[312] ^ message[315] ^ message[320] ^ message[321] ^ message[326] ^ message[328] ^ message[336] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[343] ^ message[346] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[357] ^ message[358] ^ message[361] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[369] ^ message[370] ^ message[372] ^ message[375] ^ message[377] ^ message[379] ^ message[383] ^ message[387] ^ message[388] ^ message[389] ^ message[391] ^ message[393] ^ message[394] ^ message[396] ^ message[405] ^ message[407] ^ message[409] ^ message[411] ^ message[412] ^ message[414] ^ message[417] ^ message[419] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[430] ^ message[431] ^ message[432] ^ message[433] ^ message[436] ^ message[437] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[447] ^ message[450] ^ message[451] ^ message[452] ^ message[453] ^ message[455] ^ message[456] ^ message[458] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[470] ^ message[471] ^ message[472] ^ message[476] ^ message[477] ^ message[478] ^ message[482] ^ message[490] ^ message[492] ^ message[494] ^ message[501] ^ message[504] ^ message[508] ^ message[510];
  assign _codeword[18] = message[2] ^ message[4] ^ message[9] ^ message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[22] ^ message[25] ^ message[27] ^ message[29] ^ message[31] ^ message[32] ^ message[34] ^ message[37] ^ message[38] ^ message[41] ^ message[42] ^ message[44] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[55] ^ message[60] ^ message[61] ^ message[66] ^ message[67] ^ message[69] ^ message[70] ^ message[71] ^ message[72] ^ message[76] ^ message[79] ^ message[80] ^ message[81] ^ message[83] ^ message[84] ^ message[85] ^ message[87] ^ message[89] ^ message[90] ^ message[91] ^ message[93] ^ message[95] ^ message[99] ^ message[100] ^ message[101] ^ message[104] ^ message[105] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[114] ^ message[115] ^ message[116] ^ message[119] ^ message[121] ^ message[122] ^ message[125] ^ message[126] ^ message[127] ^ message[130] ^ message[132] ^ message[134] ^ message[137] ^ message[139] ^ message[140] ^ message[141] ^ message[142] ^ message[144] ^ message[145] ^ message[146] ^ message[148] ^ message[150] ^ message[151] ^ message[152] ^ message[154] ^ message[155] ^ message[156] ^ message[158] ^ message[159] ^ message[163] ^ message[164] ^ message[167] ^ message[173] ^ message[174] ^ message[177] ^ message[178] ^ message[181] ^ message[183] ^ message[184] ^ message[187] ^ message[188] ^ message[189] ^ message[192] ^ message[195] ^ message[196] ^ message[199] ^ message[200] ^ message[202] ^ message[203] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[218] ^ message[219] ^ message[220] ^ message[223] ^ message[228] ^ message[230] ^ message[232] ^ message[233] ^ message[236] ^ message[237] ^ message[239] ^ message[240] ^ message[241] ^ message[243] ^ message[244] ^ message[250] ^ message[252] ^ message[253] ^ message[255] ^ message[256] ^ message[257] ^ message[259] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[271] ^ message[275] ^ message[278] ^ message[279] ^ message[280] ^ message[283] ^ message[289] ^ message[292] ^ message[298] ^ message[299] ^ message[302] ^ message[304] ^ message[307] ^ message[308] ^ message[311] ^ message[313] ^ message[316] ^ message[321] ^ message[322] ^ message[327] ^ message[329] ^ message[337] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[344] ^ message[347] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[358] ^ message[359] ^ message[362] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[370] ^ message[371] ^ message[373] ^ message[376] ^ message[378] ^ message[380] ^ message[384] ^ message[388] ^ message[389] ^ message[390] ^ message[392] ^ message[394] ^ message[395] ^ message[397] ^ message[406] ^ message[408] ^ message[410] ^ message[412] ^ message[413] ^ message[415] ^ message[418] ^ message[420] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[431] ^ message[432] ^ message[433] ^ message[434] ^ message[437] ^ message[438] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[448] ^ message[451] ^ message[452] ^ message[453] ^ message[454] ^ message[456] ^ message[457] ^ message[459] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[471] ^ message[472] ^ message[473] ^ message[477] ^ message[478] ^ message[479] ^ message[483] ^ message[491] ^ message[493] ^ message[495] ^ message[502] ^ message[505] ^ message[509] ^ message[511];
  assign _codeword[19] = message[0] ^ message[2] ^ message[3] ^ message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[11] ^ message[17] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[29] ^ message[30] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[51] ^ message[53] ^ message[54] ^ message[55] ^ message[56] ^ message[58] ^ message[60] ^ message[61] ^ message[63] ^ message[64] ^ message[65] ^ message[67] ^ message[68] ^ message[69] ^ message[71] ^ message[72] ^ message[79] ^ message[80] ^ message[82] ^ message[85] ^ message[91] ^ message[93] ^ message[95] ^ message[96] ^ message[97] ^ message[99] ^ message[102] ^ message[104] ^ message[105] ^ message[106] ^ message[108] ^ message[109] ^ message[111] ^ message[113] ^ message[114] ^ message[115] ^ message[122] ^ message[123] ^ message[126] ^ message[128] ^ message[131] ^ message[136] ^ message[139] ^ message[140] ^ message[143] ^ message[145] ^ message[147] ^ message[148] ^ message[150] ^ message[153] ^ message[155] ^ message[156] ^ message[157] ^ message[158] ^ message[160] ^ message[161] ^ message[163] ^ message[165] ^ message[166] ^ message[168] ^ message[169] ^ message[171] ^ message[173] ^ message[175] ^ message[176] ^ message[177] ^ message[179] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[187] ^ message[188] ^ message[191] ^ message[193] ^ message[194] ^ message[195] ^ message[197] ^ message[202] ^ message[205] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[215] ^ message[219] ^ message[220] ^ message[221] ^ message[222] ^ message[224] ^ message[226] ^ message[228] ^ message[232] ^ message[237] ^ message[238] ^ message[240] ^ message[241] ^ message[245] ^ message[246] ^ message[252] ^ message[256] ^ message[263] ^ message[266] ^ message[267] ^ message[268] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[279] ^ message[281] ^ message[282] ^ message[283] ^ message[290] ^ message[293] ^ message[294] ^ message[296] ^ message[298] ^ message[299] ^ message[302] ^ message[303] ^ message[308] ^ message[310] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[320] ^ message[321] ^ message[324] ^ message[325] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[332] ^ message[333] ^ message[334] ^ message[338] ^ message[340] ^ message[345] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[357] ^ message[358] ^ message[359] ^ message[361] ^ message[362] ^ message[365] ^ message[367] ^ message[369] ^ message[371] ^ message[372] ^ message[374] ^ message[380] ^ message[384] ^ message[386] ^ message[388] ^ message[390] ^ message[392] ^ message[395] ^ message[400] ^ message[406] ^ message[407] ^ message[408] ^ message[410] ^ message[411] ^ message[412] ^ message[415] ^ message[416] ^ message[420] ^ message[421] ^ message[423] ^ message[425] ^ message[427] ^ message[428] ^ message[430] ^ message[431] ^ message[434] ^ message[435] ^ message[439] ^ message[440] ^ message[442] ^ message[443] ^ message[445] ^ message[446] ^ message[449] ^ message[450] ^ message[451] ^ message[454] ^ message[456] ^ message[458] ^ message[459] ^ message[461] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[473] ^ message[475] ^ message[481] ^ message[484] ^ message[485] ^ message[487] ^ message[490] ^ message[495] ^ message[501] ^ message[502] ^ message[509] ^ message[510];
  assign _codeword[20] = message[1] ^ message[3] ^ message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[10] ^ message[12] ^ message[18] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[30] ^ message[31] ^ message[33] ^ message[37] ^ message[38] ^ message[41] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[52] ^ message[54] ^ message[55] ^ message[56] ^ message[57] ^ message[59] ^ message[61] ^ message[62] ^ message[64] ^ message[65] ^ message[66] ^ message[68] ^ message[69] ^ message[70] ^ message[72] ^ message[73] ^ message[80] ^ message[81] ^ message[83] ^ message[86] ^ message[92] ^ message[94] ^ message[96] ^ message[97] ^ message[98] ^ message[100] ^ message[103] ^ message[105] ^ message[106] ^ message[107] ^ message[109] ^ message[110] ^ message[112] ^ message[114] ^ message[115] ^ message[116] ^ message[123] ^ message[124] ^ message[127] ^ message[129] ^ message[132] ^ message[137] ^ message[140] ^ message[141] ^ message[144] ^ message[146] ^ message[148] ^ message[149] ^ message[151] ^ message[154] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[161] ^ message[162] ^ message[164] ^ message[166] ^ message[167] ^ message[169] ^ message[170] ^ message[172] ^ message[174] ^ message[176] ^ message[177] ^ message[178] ^ message[180] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[188] ^ message[189] ^ message[192] ^ message[194] ^ message[195] ^ message[196] ^ message[198] ^ message[203] ^ message[206] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[216] ^ message[220] ^ message[221] ^ message[222] ^ message[223] ^ message[225] ^ message[227] ^ message[229] ^ message[233] ^ message[238] ^ message[239] ^ message[241] ^ message[242] ^ message[246] ^ message[247] ^ message[253] ^ message[257] ^ message[264] ^ message[267] ^ message[268] ^ message[269] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[280] ^ message[282] ^ message[283] ^ message[284] ^ message[291] ^ message[294] ^ message[295] ^ message[297] ^ message[299] ^ message[300] ^ message[303] ^ message[304] ^ message[309] ^ message[311] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[321] ^ message[322] ^ message[325] ^ message[326] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[333] ^ message[334] ^ message[335] ^ message[339] ^ message[341] ^ message[346] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[358] ^ message[359] ^ message[360] ^ message[362] ^ message[363] ^ message[366] ^ message[368] ^ message[370] ^ message[372] ^ message[373] ^ message[375] ^ message[381] ^ message[385] ^ message[387] ^ message[389] ^ message[391] ^ message[393] ^ message[396] ^ message[401] ^ message[407] ^ message[408] ^ message[409] ^ message[411] ^ message[412] ^ message[413] ^ message[416] ^ message[417] ^ message[421] ^ message[422] ^ message[424] ^ message[426] ^ message[428] ^ message[429] ^ message[431] ^ message[432] ^ message[435] ^ message[436] ^ message[440] ^ message[441] ^ message[443] ^ message[444] ^ message[446] ^ message[447] ^ message[450] ^ message[451] ^ message[452] ^ message[455] ^ message[457] ^ message[459] ^ message[460] ^ message[462] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[474] ^ message[476] ^ message[482] ^ message[485] ^ message[486] ^ message[488] ^ message[491] ^ message[496] ^ message[502] ^ message[503] ^ message[510] ^ message[511];
  assign _codeword[21] = message[0] ^ message[5] ^ message[11] ^ message[12] ^ message[14] ^ message[17] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[40] ^ message[44] ^ message[45] ^ message[49] ^ message[50] ^ message[52] ^ message[53] ^ message[54] ^ message[56] ^ message[57] ^ message[64] ^ message[66] ^ message[67] ^ message[71] ^ message[74] ^ message[77] ^ message[79] ^ message[82] ^ message[86] ^ message[87] ^ message[88] ^ message[90] ^ message[92] ^ message[94] ^ message[98] ^ message[100] ^ message[106] ^ message[107] ^ message[109] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[120] ^ message[124] ^ message[125] ^ message[127] ^ message[128] ^ message[130] ^ message[135] ^ message[136] ^ message[139] ^ message[145] ^ message[146] ^ message[147] ^ message[148] ^ message[151] ^ message[155] ^ message[157] ^ message[160] ^ message[161] ^ message[162] ^ message[164] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[174] ^ message[175] ^ message[176] ^ message[179] ^ message[184] ^ message[186] ^ message[187] ^ message[191] ^ message[193] ^ message[194] ^ message[197] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[205] ^ message[207] ^ message[212] ^ message[213] ^ message[215] ^ message[217] ^ message[221] ^ message[223] ^ message[224] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[239] ^ message[240] ^ message[243] ^ message[244] ^ message[246] ^ message[247] ^ message[248] ^ message[251] ^ message[252] ^ message[253] ^ message[257] ^ message[260] ^ message[264] ^ message[268] ^ message[270] ^ message[272] ^ message[273] ^ message[274] ^ message[276] ^ message[277] ^ message[278] ^ message[280] ^ message[281] ^ message[282] ^ message[285] ^ message[292] ^ message[294] ^ message[295] ^ message[301] ^ message[302] ^ message[304] ^ message[309] ^ message[312] ^ message[313] ^ message[314] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[324] ^ message[325] ^ message[326] ^ message[330] ^ message[331] ^ message[333] ^ message[335] ^ message[336] ^ message[340] ^ message[341] ^ message[343] ^ message[347] ^ message[348] ^ message[350] ^ message[352] ^ message[353] ^ message[354] ^ message[357] ^ message[358] ^ message[359] ^ message[362] ^ message[364] ^ message[366] ^ message[367] ^ message[368] ^ message[371] ^ message[373] ^ message[374] ^ message[376] ^ message[377] ^ message[379] ^ message[380] ^ message[381] ^ message[382] ^ message[384] ^ message[385] ^ message[389] ^ message[390] ^ message[391] ^ message[393] ^ message[394] ^ message[396] ^ message[397] ^ message[398] ^ message[400] ^ message[402] ^ message[406] ^ message[415] ^ message[417] ^ message[418] ^ message[419] ^ message[420] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[430] ^ message[431] ^ message[436] ^ message[437] ^ message[438] ^ message[440] ^ message[441] ^ message[445] ^ message[447] ^ message[448] ^ message[450] ^ message[455] ^ message[457] ^ message[458] ^ message[459] ^ message[463] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[472] ^ message[474] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[483] ^ message[485] ^ message[486] ^ message[489] ^ message[490] ^ message[494] ^ message[495] ^ message[496] ^ message[497] ^ message[501] ^ message[502] ^ message[504] ^ message[506] ^ message[509] ^ message[511];
  assign _codeword[22] = message[1] ^ message[6] ^ message[12] ^ message[13] ^ message[15] ^ message[18] ^ message[20] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[32] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[41] ^ message[45] ^ message[46] ^ message[50] ^ message[51] ^ message[53] ^ message[54] ^ message[55] ^ message[57] ^ message[58] ^ message[65] ^ message[67] ^ message[68] ^ message[72] ^ message[75] ^ message[78] ^ message[80] ^ message[83] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[93] ^ message[95] ^ message[99] ^ message[101] ^ message[107] ^ message[108] ^ message[110] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[121] ^ message[125] ^ message[126] ^ message[128] ^ message[129] ^ message[131] ^ message[136] ^ message[137] ^ message[140] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[152] ^ message[156] ^ message[158] ^ message[161] ^ message[162] ^ message[163] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[175] ^ message[176] ^ message[177] ^ message[180] ^ message[185] ^ message[187] ^ message[188] ^ message[192] ^ message[194] ^ message[195] ^ message[198] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[206] ^ message[208] ^ message[213] ^ message[214] ^ message[216] ^ message[218] ^ message[222] ^ message[224] ^ message[225] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[240] ^ message[241] ^ message[244] ^ message[245] ^ message[247] ^ message[248] ^ message[249] ^ message[252] ^ message[253] ^ message[254] ^ message[258] ^ message[261] ^ message[265] ^ message[269] ^ message[271] ^ message[273] ^ message[274] ^ message[275] ^ message[277] ^ message[278] ^ message[279] ^ message[281] ^ message[282] ^ message[283] ^ message[286] ^ message[293] ^ message[295] ^ message[296] ^ message[302] ^ message[303] ^ message[305] ^ message[310] ^ message[313] ^ message[314] ^ message[315] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[325] ^ message[326] ^ message[327] ^ message[331] ^ message[332] ^ message[334] ^ message[336] ^ message[337] ^ message[341] ^ message[342] ^ message[344] ^ message[348] ^ message[349] ^ message[351] ^ message[353] ^ message[354] ^ message[355] ^ message[358] ^ message[359] ^ message[360] ^ message[363] ^ message[365] ^ message[367] ^ message[368] ^ message[369] ^ message[372] ^ message[374] ^ message[375] ^ message[377] ^ message[378] ^ message[380] ^ message[381] ^ message[382] ^ message[383] ^ message[385] ^ message[386] ^ message[390] ^ message[391] ^ message[392] ^ message[394] ^ message[395] ^ message[397] ^ message[398] ^ message[399] ^ message[401] ^ message[403] ^ message[407] ^ message[416] ^ message[418] ^ message[419] ^ message[420] ^ message[421] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[431] ^ message[432] ^ message[437] ^ message[438] ^ message[439] ^ message[441] ^ message[442] ^ message[446] ^ message[448] ^ message[449] ^ message[451] ^ message[456] ^ message[458] ^ message[459] ^ message[460] ^ message[464] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[473] ^ message[475] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[484] ^ message[486] ^ message[487] ^ message[490] ^ message[491] ^ message[495] ^ message[496] ^ message[497] ^ message[498] ^ message[502] ^ message[503] ^ message[505] ^ message[507] ^ message[510];
  assign _codeword[23] = message[0] ^ message[4] ^ message[6] ^ message[8] ^ message[9] ^ message[10] ^ message[12] ^ message[16] ^ message[17] ^ message[19] ^ message[21] ^ message[23] ^ message[24] ^ message[26] ^ message[29] ^ message[34] ^ message[40] ^ message[44] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[56] ^ message[59] ^ message[60] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[68] ^ message[70] ^ message[76] ^ message[77] ^ message[86] ^ message[89] ^ message[93] ^ message[95] ^ message[96] ^ message[97] ^ message[99] ^ message[101] ^ message[102] ^ message[104] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[115] ^ message[120] ^ message[122] ^ message[126] ^ message[129] ^ message[130] ^ message[132] ^ message[133] ^ message[135] ^ message[136] ^ message[137] ^ message[139] ^ message[142] ^ message[146] ^ message[147] ^ message[151] ^ message[152] ^ message[153] ^ message[157] ^ message[158] ^ message[161] ^ message[162] ^ message[167] ^ message[168] ^ message[170] ^ message[172] ^ message[173] ^ message[174] ^ message[183] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[190] ^ message[191] ^ message[193] ^ message[194] ^ message[199] ^ message[200] ^ message[207] ^ message[209] ^ message[215] ^ message[217] ^ message[219] ^ message[222] ^ message[223] ^ message[225] ^ message[228] ^ message[229] ^ message[235] ^ message[241] ^ message[244] ^ message[245] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[255] ^ message[257] ^ message[258] ^ message[259] ^ message[260] ^ message[262] ^ message[264] ^ message[265] ^ message[266] ^ message[269] ^ message[270] ^ message[273] ^ message[276] ^ message[278] ^ message[279] ^ message[287] ^ message[297] ^ message[298] ^ message[300] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[309] ^ message[310] ^ message[311] ^ message[313] ^ message[314] ^ message[319] ^ message[324] ^ message[325] ^ message[326] ^ message[328] ^ message[329] ^ message[334] ^ message[335] ^ message[337] ^ message[338] ^ message[341] ^ message[345] ^ message[348] ^ message[349] ^ message[352] ^ message[354] ^ message[357] ^ message[358] ^ message[359] ^ message[362] ^ message[363] ^ message[364] ^ message[370] ^ message[373] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[380] ^ message[382] ^ message[383] ^ message[385] ^ message[387] ^ message[388] ^ message[389] ^ message[395] ^ message[399] ^ message[402] ^ message[404] ^ message[406] ^ message[409] ^ message[410] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[417] ^ message[421] ^ message[422] ^ message[425] ^ message[427] ^ message[428] ^ message[431] ^ message[439] ^ message[443] ^ message[444] ^ message[447] ^ message[449] ^ message[451] ^ message[453] ^ message[455] ^ message[456] ^ message[465] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[472] ^ message[475] ^ message[476] ^ message[478] ^ message[482] ^ message[483] ^ message[488] ^ message[490] ^ message[491] ^ message[494] ^ message[495] ^ message[497] ^ message[498] ^ message[499] ^ message[501] ^ message[502] ^ message[504] ^ message[508] ^ message[509] ^ message[511];
  assign _codeword[24] = message[1] ^ message[5] ^ message[7] ^ message[9] ^ message[10] ^ message[11] ^ message[13] ^ message[17] ^ message[18] ^ message[20] ^ message[22] ^ message[24] ^ message[25] ^ message[27] ^ message[30] ^ message[35] ^ message[41] ^ message[45] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[57] ^ message[60] ^ message[61] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[69] ^ message[71] ^ message[77] ^ message[78] ^ message[87] ^ message[90] ^ message[94] ^ message[96] ^ message[97] ^ message[98] ^ message[100] ^ message[102] ^ message[103] ^ message[105] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[116] ^ message[121] ^ message[123] ^ message[127] ^ message[130] ^ message[131] ^ message[133] ^ message[134] ^ message[136] ^ message[137] ^ message[138] ^ message[140] ^ message[143] ^ message[147] ^ message[148] ^ message[152] ^ message[153] ^ message[154] ^ message[158] ^ message[159] ^ message[162] ^ message[163] ^ message[168] ^ message[169] ^ message[171] ^ message[173] ^ message[174] ^ message[175] ^ message[184] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[200] ^ message[201] ^ message[208] ^ message[210] ^ message[216] ^ message[218] ^ message[220] ^ message[223] ^ message[224] ^ message[226] ^ message[229] ^ message[230] ^ message[236] ^ message[242] ^ message[245] ^ message[246] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[256] ^ message[258] ^ message[259] ^ message[260] ^ message[261] ^ message[263] ^ message[265] ^ message[266] ^ message[267] ^ message[270] ^ message[271] ^ message[274] ^ message[277] ^ message[279] ^ message[280] ^ message[288] ^ message[298] ^ message[299] ^ message[301] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[310] ^ message[311] ^ message[312] ^ message[314] ^ message[315] ^ message[320] ^ message[325] ^ message[326] ^ message[327] ^ message[329] ^ message[330] ^ message[335] ^ message[336] ^ message[338] ^ message[339] ^ message[342] ^ message[346] ^ message[349] ^ message[350] ^ message[353] ^ message[355] ^ message[358] ^ message[359] ^ message[360] ^ message[363] ^ message[364] ^ message[365] ^ message[371] ^ message[374] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[381] ^ message[383] ^ message[384] ^ message[386] ^ message[388] ^ message[389] ^ message[390] ^ message[396] ^ message[400] ^ message[403] ^ message[405] ^ message[407] ^ message[410] ^ message[411] ^ message[413] ^ message[414] ^ message[415] ^ message[416] ^ message[418] ^ message[422] ^ message[423] ^ message[426] ^ message[428] ^ message[429] ^ message[432] ^ message[440] ^ message[444] ^ message[445] ^ message[448] ^ message[450] ^ message[452] ^ message[454] ^ message[456] ^ message[457] ^ message[466] ^ message[469] ^ message[470] ^ message[471] ^ message[472] ^ message[473] ^ message[476] ^ message[477] ^ message[479] ^ message[483] ^ message[484] ^ message[489] ^ message[491] ^ message[492] ^ message[495] ^ message[496] ^ message[498] ^ message[499] ^ message[500] ^ message[502] ^ message[503] ^ message[505] ^ message[509] ^ message[510];
  assign _codeword[25] = message[2] ^ message[6] ^ message[8] ^ message[10] ^ message[11] ^ message[12] ^ message[14] ^ message[18] ^ message[19] ^ message[21] ^ message[23] ^ message[25] ^ message[26] ^ message[28] ^ message[31] ^ message[36] ^ message[42] ^ message[46] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[58] ^ message[61] ^ message[62] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[70] ^ message[72] ^ message[78] ^ message[79] ^ message[88] ^ message[91] ^ message[95] ^ message[97] ^ message[98] ^ message[99] ^ message[101] ^ message[103] ^ message[104] ^ message[106] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[117] ^ message[122] ^ message[124] ^ message[128] ^ message[131] ^ message[132] ^ message[134] ^ message[135] ^ message[137] ^ message[138] ^ message[139] ^ message[141] ^ message[144] ^ message[148] ^ message[149] ^ message[153] ^ message[154] ^ message[155] ^ message[159] ^ message[160] ^ message[163] ^ message[164] ^ message[169] ^ message[170] ^ message[172] ^ message[174] ^ message[175] ^ message[176] ^ message[185] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[192] ^ message[193] ^ message[195] ^ message[196] ^ message[201] ^ message[202] ^ message[209] ^ message[211] ^ message[217] ^ message[219] ^ message[221] ^ message[224] ^ message[225] ^ message[227] ^ message[230] ^ message[231] ^ message[237] ^ message[243] ^ message[246] ^ message[247] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[257] ^ message[259] ^ message[260] ^ message[261] ^ message[262] ^ message[264] ^ message[266] ^ message[267] ^ message[268] ^ message[271] ^ message[272] ^ message[275] ^ message[278] ^ message[280] ^ message[281] ^ message[289] ^ message[299] ^ message[300] ^ message[302] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[311] ^ message[312] ^ message[313] ^ message[315] ^ message[316] ^ message[321] ^ message[326] ^ message[327] ^ message[328] ^ message[330] ^ message[331] ^ message[336] ^ message[337] ^ message[339] ^ message[340] ^ message[343] ^ message[347] ^ message[350] ^ message[351] ^ message[354] ^ message[356] ^ message[359] ^ message[360] ^ message[361] ^ message[364] ^ message[365] ^ message[366] ^ message[372] ^ message[375] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[382] ^ message[384] ^ message[385] ^ message[387] ^ message[389] ^ message[390] ^ message[391] ^ message[397] ^ message[401] ^ message[404] ^ message[406] ^ message[408] ^ message[411] ^ message[412] ^ message[414] ^ message[415] ^ message[416] ^ message[417] ^ message[419] ^ message[423] ^ message[424] ^ message[427] ^ message[429] ^ message[430] ^ message[433] ^ message[441] ^ message[445] ^ message[446] ^ message[449] ^ message[451] ^ message[453] ^ message[455] ^ message[457] ^ message[458] ^ message[467] ^ message[470] ^ message[471] ^ message[472] ^ message[473] ^ message[474] ^ message[477] ^ message[478] ^ message[480] ^ message[484] ^ message[485] ^ message[490] ^ message[492] ^ message[493] ^ message[496] ^ message[497] ^ message[499] ^ message[500] ^ message[501] ^ message[503] ^ message[504] ^ message[506] ^ message[510] ^ message[511];
  assign _codeword[26] = message[3] ^ message[7] ^ message[9] ^ message[11] ^ message[12] ^ message[13] ^ message[15] ^ message[19] ^ message[20] ^ message[22] ^ message[24] ^ message[26] ^ message[27] ^ message[29] ^ message[32] ^ message[37] ^ message[43] ^ message[47] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[59] ^ message[62] ^ message[63] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[71] ^ message[73] ^ message[79] ^ message[80] ^ message[89] ^ message[92] ^ message[96] ^ message[98] ^ message[99] ^ message[100] ^ message[102] ^ message[104] ^ message[105] ^ message[107] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[118] ^ message[123] ^ message[125] ^ message[129] ^ message[132] ^ message[133] ^ message[135] ^ message[136] ^ message[138] ^ message[139] ^ message[140] ^ message[142] ^ message[145] ^ message[149] ^ message[150] ^ message[154] ^ message[155] ^ message[156] ^ message[160] ^ message[161] ^ message[164] ^ message[165] ^ message[170] ^ message[171] ^ message[173] ^ message[175] ^ message[176] ^ message[177] ^ message[186] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[193] ^ message[194] ^ message[196] ^ message[197] ^ message[202] ^ message[203] ^ message[210] ^ message[212] ^ message[218] ^ message[220] ^ message[222] ^ message[225] ^ message[226] ^ message[228] ^ message[231] ^ message[232] ^ message[238] ^ message[244] ^ message[247] ^ message[248] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[258] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[265] ^ message[267] ^ message[268] ^ message[269] ^ message[272] ^ message[273] ^ message[276] ^ message[279] ^ message[281] ^ message[282] ^ message[290] ^ message[300] ^ message[301] ^ message[303] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[312] ^ message[313] ^ message[314] ^ message[316] ^ message[317] ^ message[322] ^ message[327] ^ message[328] ^ message[329] ^ message[331] ^ message[332] ^ message[337] ^ message[338] ^ message[340] ^ message[341] ^ message[344] ^ message[348] ^ message[351] ^ message[352] ^ message[355] ^ message[357] ^ message[360] ^ message[361] ^ message[362] ^ message[365] ^ message[366] ^ message[367] ^ message[373] ^ message[376] ^ message[378] ^ message[379] ^ message[380] ^ message[381] ^ message[383] ^ message[385] ^ message[386] ^ message[388] ^ message[390] ^ message[391] ^ message[392] ^ message[398] ^ message[402] ^ message[405] ^ message[407] ^ message[409] ^ message[412] ^ message[413] ^ message[415] ^ message[416] ^ message[417] ^ message[418] ^ message[420] ^ message[424] ^ message[425] ^ message[428] ^ message[430] ^ message[431] ^ message[434] ^ message[442] ^ message[446] ^ message[447] ^ message[450] ^ message[452] ^ message[454] ^ message[456] ^ message[458] ^ message[459] ^ message[468] ^ message[471] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[478] ^ message[479] ^ message[481] ^ message[485] ^ message[486] ^ message[491] ^ message[493] ^ message[494] ^ message[497] ^ message[498] ^ message[500] ^ message[501] ^ message[502] ^ message[504] ^ message[505] ^ message[507] ^ message[511];
  assign _codeword[27] = message[4] ^ message[8] ^ message[10] ^ message[12] ^ message[13] ^ message[14] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[25] ^ message[27] ^ message[28] ^ message[30] ^ message[33] ^ message[38] ^ message[44] ^ message[48] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[60] ^ message[63] ^ message[64] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[72] ^ message[74] ^ message[80] ^ message[81] ^ message[90] ^ message[93] ^ message[97] ^ message[99] ^ message[100] ^ message[101] ^ message[103] ^ message[105] ^ message[106] ^ message[108] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[119] ^ message[124] ^ message[126] ^ message[130] ^ message[133] ^ message[134] ^ message[136] ^ message[137] ^ message[139] ^ message[140] ^ message[141] ^ message[143] ^ message[146] ^ message[150] ^ message[151] ^ message[155] ^ message[156] ^ message[157] ^ message[161] ^ message[162] ^ message[165] ^ message[166] ^ message[171] ^ message[172] ^ message[174] ^ message[176] ^ message[177] ^ message[178] ^ message[187] ^ message[189] ^ message[190] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[197] ^ message[198] ^ message[203] ^ message[204] ^ message[211] ^ message[213] ^ message[219] ^ message[221] ^ message[223] ^ message[226] ^ message[227] ^ message[229] ^ message[232] ^ message[233] ^ message[239] ^ message[245] ^ message[248] ^ message[249] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[256] ^ message[259] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[266] ^ message[268] ^ message[269] ^ message[270] ^ message[273] ^ message[274] ^ message[277] ^ message[280] ^ message[282] ^ message[283] ^ message[291] ^ message[301] ^ message[302] ^ message[304] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[313] ^ message[314] ^ message[315] ^ message[317] ^ message[318] ^ message[323] ^ message[328] ^ message[329] ^ message[330] ^ message[332] ^ message[333] ^ message[338] ^ message[339] ^ message[341] ^ message[342] ^ message[345] ^ message[349] ^ message[352] ^ message[353] ^ message[356] ^ message[358] ^ message[361] ^ message[362] ^ message[363] ^ message[366] ^ message[367] ^ message[368] ^ message[374] ^ message[377] ^ message[379] ^ message[380] ^ message[381] ^ message[382] ^ message[384] ^ message[386] ^ message[387] ^ message[389] ^ message[391] ^ message[392] ^ message[393] ^ message[399] ^ message[403] ^ message[406] ^ message[408] ^ message[410] ^ message[413] ^ message[414] ^ message[416] ^ message[417] ^ message[418] ^ message[419] ^ message[421] ^ message[425] ^ message[426] ^ message[429] ^ message[431] ^ message[432] ^ message[435] ^ message[443] ^ message[447] ^ message[448] ^ message[451] ^ message[453] ^ message[455] ^ message[457] ^ message[459] ^ message[460] ^ message[469] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[479] ^ message[480] ^ message[482] ^ message[486] ^ message[487] ^ message[492] ^ message[494] ^ message[495] ^ message[498] ^ message[499] ^ message[501] ^ message[502] ^ message[503] ^ message[505] ^ message[506] ^ message[508];
  assign _codeword[28] = message[0] ^ message[2] ^ message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[10] ^ message[11] ^ message[12] ^ message[15] ^ message[21] ^ message[22] ^ message[23] ^ message[25] ^ message[26] ^ message[27] ^ message[31] ^ message[33] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[40] ^ message[42] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[50] ^ message[52] ^ message[53] ^ message[56] ^ message[58] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[67] ^ message[68] ^ message[71] ^ message[75] ^ message[77] ^ message[79] ^ message[82] ^ message[84] ^ message[86] ^ message[88] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[95] ^ message[97] ^ message[98] ^ message[99] ^ message[102] ^ message[106] ^ message[107] ^ message[108] ^ message[110] ^ message[112] ^ message[114] ^ message[115] ^ message[118] ^ message[125] ^ message[131] ^ message[133] ^ message[134] ^ message[136] ^ message[137] ^ message[139] ^ message[140] ^ message[144] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[156] ^ message[157] ^ message[159] ^ message[161] ^ message[162] ^ message[164] ^ message[167] ^ message[169] ^ message[171] ^ message[172] ^ message[174] ^ message[175] ^ message[176] ^ message[179] ^ message[181] ^ message[183] ^ message[185] ^ message[187] ^ message[188] ^ message[189] ^ message[192] ^ message[193] ^ message[194] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[212] ^ message[220] ^ message[224] ^ message[226] ^ message[227] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[240] ^ message[242] ^ message[244] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[255] ^ message[256] ^ message[258] ^ message[262] ^ message[263] ^ message[267] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[278] ^ message[280] ^ message[281] ^ message[282] ^ message[292] ^ message[294] ^ message[296] ^ message[298] ^ message[300] ^ message[303] ^ message[307] ^ message[308] ^ message[311] ^ message[313] ^ message[314] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[325] ^ message[327] ^ message[330] ^ message[331] ^ message[332] ^ message[339] ^ message[340] ^ message[341] ^ message[346] ^ message[348] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[358] ^ message[359] ^ message[360] ^ message[361] ^ message[364] ^ message[366] ^ message[367] ^ message[375] ^ message[377] ^ message[378] ^ message[379] ^ message[382] ^ message[383] ^ message[384] ^ message[386] ^ message[387] ^ message[389] ^ message[390] ^ message[391] ^ message[394] ^ message[396] ^ message[398] ^ message[404] ^ message[406] ^ message[407] ^ message[408] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[417] ^ message[418] ^ message[422] ^ message[424] ^ message[427] ^ message[429] ^ message[430] ^ message[431] ^ message[436] ^ message[438] ^ message[440] ^ message[442] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[453] ^ message[454] ^ message[455] ^ message[457] ^ message[458] ^ message[459] ^ message[470] ^ message[472] ^ message[473] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[483] ^ message[485] ^ message[488] ^ message[490] ^ message[492] ^ message[493] ^ message[494] ^ message[499] ^ message[500] ^ message[501] ^ message[504] ^ message[507];
  assign _codeword[29] = message[1] ^ message[3] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[11] ^ message[12] ^ message[13] ^ message[16] ^ message[22] ^ message[23] ^ message[24] ^ message[26] ^ message[27] ^ message[28] ^ message[32] ^ message[34] ^ message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[41] ^ message[43] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[51] ^ message[53] ^ message[54] ^ message[57] ^ message[59] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[68] ^ message[69] ^ message[72] ^ message[76] ^ message[78] ^ message[80] ^ message[83] ^ message[85] ^ message[87] ^ message[89] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[96] ^ message[98] ^ message[99] ^ message[100] ^ message[103] ^ message[107] ^ message[108] ^ message[109] ^ message[111] ^ message[113] ^ message[115] ^ message[116] ^ message[119] ^ message[126] ^ message[132] ^ message[134] ^ message[135] ^ message[137] ^ message[138] ^ message[140] ^ message[141] ^ message[145] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[157] ^ message[158] ^ message[160] ^ message[162] ^ message[163] ^ message[165] ^ message[168] ^ message[170] ^ message[172] ^ message[173] ^ message[175] ^ message[176] ^ message[177] ^ message[180] ^ message[182] ^ message[184] ^ message[186] ^ message[188] ^ message[189] ^ message[190] ^ message[193] ^ message[194] ^ message[195] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[213] ^ message[221] ^ message[225] ^ message[227] ^ message[228] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[241] ^ message[243] ^ message[245] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[256] ^ message[257] ^ message[259] ^ message[263] ^ message[264] ^ message[268] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[279] ^ message[281] ^ message[282] ^ message[283] ^ message[293] ^ message[295] ^ message[297] ^ message[299] ^ message[301] ^ message[304] ^ message[308] ^ message[309] ^ message[312] ^ message[314] ^ message[315] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[326] ^ message[328] ^ message[331] ^ message[332] ^ message[333] ^ message[340] ^ message[341] ^ message[342] ^ message[347] ^ message[349] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[359] ^ message[360] ^ message[361] ^ message[362] ^ message[365] ^ message[367] ^ message[368] ^ message[376] ^ message[378] ^ message[379] ^ message[380] ^ message[383] ^ message[384] ^ message[385] ^ message[387] ^ message[388] ^ message[390] ^ message[391] ^ message[392] ^ message[395] ^ message[397] ^ message[399] ^ message[405] ^ message[407] ^ message[408] ^ message[409] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[418] ^ message[419] ^ message[423] ^ message[425] ^ message[428] ^ message[430] ^ message[431] ^ message[432] ^ message[437] ^ message[439] ^ message[441] ^ message[443] ^ message[449] ^ message[450] ^ message[451] ^ message[452] ^ message[454] ^ message[455] ^ message[456] ^ message[458] ^ message[459] ^ message[460] ^ message[471] ^ message[473] ^ message[474] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[484] ^ message[486] ^ message[489] ^ message[491] ^ message[493] ^ message[494] ^ message[495] ^ message[500] ^ message[501] ^ message[502] ^ message[505] ^ message[508];
  assign _codeword[30] = message[0];
  assign _codeword[31] = message[1];
  assign _codeword[32] = message[2];
  assign _codeword[33] = message[3];
  assign _codeword[34] = message[4];
  assign _codeword[35] = message[5];
  assign _codeword[36] = message[6];
  assign _codeword[37] = message[7];
  assign _codeword[38] = message[8];
  assign _codeword[39] = message[9];
  assign _codeword[40] = message[10];
  assign _codeword[41] = message[11];
  assign _codeword[42] = message[12];
  assign _codeword[43] = message[13];
  assign _codeword[44] = message[14];
  assign _codeword[45] = message[15];
  assign _codeword[46] = message[16];
  assign _codeword[47] = message[17];
  assign _codeword[48] = message[18];
  assign _codeword[49] = message[19];
  assign _codeword[50] = message[20];
  assign _codeword[51] = message[21];
  assign _codeword[52] = message[22];
  assign _codeword[53] = message[23];
  assign _codeword[54] = message[24];
  assign _codeword[55] = message[25];
  assign _codeword[56] = message[26];
  assign _codeword[57] = message[27];
  assign _codeword[58] = message[28];
  assign _codeword[59] = message[29];
  assign _codeword[60] = message[30];
  assign _codeword[61] = message[31];
  assign _codeword[62] = message[32];
  assign _codeword[63] = message[33];
  assign _codeword[64] = message[34];
  assign _codeword[65] = message[35];
  assign _codeword[66] = message[36];
  assign _codeword[67] = message[37];
  assign _codeword[68] = message[38];
  assign _codeword[69] = message[39];
  assign _codeword[70] = message[40];
  assign _codeword[71] = message[41];
  assign _codeword[72] = message[42];
  assign _codeword[73] = message[43];
  assign _codeword[74] = message[44];
  assign _codeword[75] = message[45];
  assign _codeword[76] = message[46];
  assign _codeword[77] = message[47];
  assign _codeword[78] = message[48];
  assign _codeword[79] = message[49];
  assign _codeword[80] = message[50];
  assign _codeword[81] = message[51];
  assign _codeword[82] = message[52];
  assign _codeword[83] = message[53];
  assign _codeword[84] = message[54];
  assign _codeword[85] = message[55];
  assign _codeword[86] = message[56];
  assign _codeword[87] = message[57];
  assign _codeword[88] = message[58];
  assign _codeword[89] = message[59];
  assign _codeword[90] = message[60];
  assign _codeword[91] = message[61];
  assign _codeword[92] = message[62];
  assign _codeword[93] = message[63];
  assign _codeword[94] = message[64];
  assign _codeword[95] = message[65];
  assign _codeword[96] = message[66];
  assign _codeword[97] = message[67];
  assign _codeword[98] = message[68];
  assign _codeword[99] = message[69];
  assign _codeword[100] = message[70];
  assign _codeword[101] = message[71];
  assign _codeword[102] = message[72];
  assign _codeword[103] = message[73];
  assign _codeword[104] = message[74];
  assign _codeword[105] = message[75];
  assign _codeword[106] = message[76];
  assign _codeword[107] = message[77];
  assign _codeword[108] = message[78];
  assign _codeword[109] = message[79];
  assign _codeword[110] = message[80];
  assign _codeword[111] = message[81];
  assign _codeword[112] = message[82];
  assign _codeword[113] = message[83];
  assign _codeword[114] = message[84];
  assign _codeword[115] = message[85];
  assign _codeword[116] = message[86];
  assign _codeword[117] = message[87];
  assign _codeword[118] = message[88];
  assign _codeword[119] = message[89];
  assign _codeword[120] = message[90];
  assign _codeword[121] = message[91];
  assign _codeword[122] = message[92];
  assign _codeword[123] = message[93];
  assign _codeword[124] = message[94];
  assign _codeword[125] = message[95];
  assign _codeword[126] = message[96];
  assign _codeword[127] = message[97];
  assign _codeword[128] = message[98];
  assign _codeword[129] = message[99];
  assign _codeword[130] = message[100];
  assign _codeword[131] = message[101];
  assign _codeword[132] = message[102];
  assign _codeword[133] = message[103];
  assign _codeword[134] = message[104];
  assign _codeword[135] = message[105];
  assign _codeword[136] = message[106];
  assign _codeword[137] = message[107];
  assign _codeword[138] = message[108];
  assign _codeword[139] = message[109];
  assign _codeword[140] = message[110];
  assign _codeword[141] = message[111];
  assign _codeword[142] = message[112];
  assign _codeword[143] = message[113];
  assign _codeword[144] = message[114];
  assign _codeword[145] = message[115];
  assign _codeword[146] = message[116];
  assign _codeword[147] = message[117];
  assign _codeword[148] = message[118];
  assign _codeword[149] = message[119];
  assign _codeword[150] = message[120];
  assign _codeword[151] = message[121];
  assign _codeword[152] = message[122];
  assign _codeword[153] = message[123];
  assign _codeword[154] = message[124];
  assign _codeword[155] = message[125];
  assign _codeword[156] = message[126];
  assign _codeword[157] = message[127];
  assign _codeword[158] = message[128];
  assign _codeword[159] = message[129];
  assign _codeword[160] = message[130];
  assign _codeword[161] = message[131];
  assign _codeword[162] = message[132];
  assign _codeword[163] = message[133];
  assign _codeword[164] = message[134];
  assign _codeword[165] = message[135];
  assign _codeword[166] = message[136];
  assign _codeword[167] = message[137];
  assign _codeword[168] = message[138];
  assign _codeword[169] = message[139];
  assign _codeword[170] = message[140];
  assign _codeword[171] = message[141];
  assign _codeword[172] = message[142];
  assign _codeword[173] = message[143];
  assign _codeword[174] = message[144];
  assign _codeword[175] = message[145];
  assign _codeword[176] = message[146];
  assign _codeword[177] = message[147];
  assign _codeword[178] = message[148];
  assign _codeword[179] = message[149];
  assign _codeword[180] = message[150];
  assign _codeword[181] = message[151];
  assign _codeword[182] = message[152];
  assign _codeword[183] = message[153];
  assign _codeword[184] = message[154];
  assign _codeword[185] = message[155];
  assign _codeword[186] = message[156];
  assign _codeword[187] = message[157];
  assign _codeword[188] = message[158];
  assign _codeword[189] = message[159];
  assign _codeword[190] = message[160];
  assign _codeword[191] = message[161];
  assign _codeword[192] = message[162];
  assign _codeword[193] = message[163];
  assign _codeword[194] = message[164];
  assign _codeword[195] = message[165];
  assign _codeword[196] = message[166];
  assign _codeword[197] = message[167];
  assign _codeword[198] = message[168];
  assign _codeword[199] = message[169];
  assign _codeword[200] = message[170];
  assign _codeword[201] = message[171];
  assign _codeword[202] = message[172];
  assign _codeword[203] = message[173];
  assign _codeword[204] = message[174];
  assign _codeword[205] = message[175];
  assign _codeword[206] = message[176];
  assign _codeword[207] = message[177];
  assign _codeword[208] = message[178];
  assign _codeword[209] = message[179];
  assign _codeword[210] = message[180];
  assign _codeword[211] = message[181];
  assign _codeword[212] = message[182];
  assign _codeword[213] = message[183];
  assign _codeword[214] = message[184];
  assign _codeword[215] = message[185];
  assign _codeword[216] = message[186];
  assign _codeword[217] = message[187];
  assign _codeword[218] = message[188];
  assign _codeword[219] = message[189];
  assign _codeword[220] = message[190];
  assign _codeword[221] = message[191];
  assign _codeword[222] = message[192];
  assign _codeword[223] = message[193];
  assign _codeword[224] = message[194];
  assign _codeword[225] = message[195];
  assign _codeword[226] = message[196];
  assign _codeword[227] = message[197];
  assign _codeword[228] = message[198];
  assign _codeword[229] = message[199];
  assign _codeword[230] = message[200];
  assign _codeword[231] = message[201];
  assign _codeword[232] = message[202];
  assign _codeword[233] = message[203];
  assign _codeword[234] = message[204];
  assign _codeword[235] = message[205];
  assign _codeword[236] = message[206];
  assign _codeword[237] = message[207];
  assign _codeword[238] = message[208];
  assign _codeword[239] = message[209];
  assign _codeword[240] = message[210];
  assign _codeword[241] = message[211];
  assign _codeword[242] = message[212];
  assign _codeword[243] = message[213];
  assign _codeword[244] = message[214];
  assign _codeword[245] = message[215];
  assign _codeword[246] = message[216];
  assign _codeword[247] = message[217];
  assign _codeword[248] = message[218];
  assign _codeword[249] = message[219];
  assign _codeword[250] = message[220];
  assign _codeword[251] = message[221];
  assign _codeword[252] = message[222];
  assign _codeword[253] = message[223];
  assign _codeword[254] = message[224];
  assign _codeword[255] = message[225];
  assign _codeword[256] = message[226];
  assign _codeword[257] = message[227];
  assign _codeword[258] = message[228];
  assign _codeword[259] = message[229];
  assign _codeword[260] = message[230];
  assign _codeword[261] = message[231];
  assign _codeword[262] = message[232];
  assign _codeword[263] = message[233];
  assign _codeword[264] = message[234];
  assign _codeword[265] = message[235];
  assign _codeword[266] = message[236];
  assign _codeword[267] = message[237];
  assign _codeword[268] = message[238];
  assign _codeword[269] = message[239];
  assign _codeword[270] = message[240];
  assign _codeword[271] = message[241];
  assign _codeword[272] = message[242];
  assign _codeword[273] = message[243];
  assign _codeword[274] = message[244];
  assign _codeword[275] = message[245];
  assign _codeword[276] = message[246];
  assign _codeword[277] = message[247];
  assign _codeword[278] = message[248];
  assign _codeword[279] = message[249];
  assign _codeword[280] = message[250];
  assign _codeword[281] = message[251];
  assign _codeword[282] = message[252];
  assign _codeword[283] = message[253];
  assign _codeword[284] = message[254];
  assign _codeword[285] = message[255];
  assign _codeword[286] = message[256];
  assign _codeword[287] = message[257];
  assign _codeword[288] = message[258];
  assign _codeword[289] = message[259];
  assign _codeword[290] = message[260];
  assign _codeword[291] = message[261];
  assign _codeword[292] = message[262];
  assign _codeword[293] = message[263];
  assign _codeword[294] = message[264];
  assign _codeword[295] = message[265];
  assign _codeword[296] = message[266];
  assign _codeword[297] = message[267];
  assign _codeword[298] = message[268];
  assign _codeword[299] = message[269];
  assign _codeword[300] = message[270];
  assign _codeword[301] = message[271];
  assign _codeword[302] = message[272];
  assign _codeword[303] = message[273];
  assign _codeword[304] = message[274];
  assign _codeword[305] = message[275];
  assign _codeword[306] = message[276];
  assign _codeword[307] = message[277];
  assign _codeword[308] = message[278];
  assign _codeword[309] = message[279];
  assign _codeword[310] = message[280];
  assign _codeword[311] = message[281];
  assign _codeword[312] = message[282];
  assign _codeword[313] = message[283];
  assign _codeword[314] = message[284];
  assign _codeword[315] = message[285];
  assign _codeword[316] = message[286];
  assign _codeword[317] = message[287];
  assign _codeword[318] = message[288];
  assign _codeword[319] = message[289];
  assign _codeword[320] = message[290];
  assign _codeword[321] = message[291];
  assign _codeword[322] = message[292];
  assign _codeword[323] = message[293];
  assign _codeword[324] = message[294];
  assign _codeword[325] = message[295];
  assign _codeword[326] = message[296];
  assign _codeword[327] = message[297];
  assign _codeword[328] = message[298];
  assign _codeword[329] = message[299];
  assign _codeword[330] = message[300];
  assign _codeword[331] = message[301];
  assign _codeword[332] = message[302];
  assign _codeword[333] = message[303];
  assign _codeword[334] = message[304];
  assign _codeword[335] = message[305];
  assign _codeword[336] = message[306];
  assign _codeword[337] = message[307];
  assign _codeword[338] = message[308];
  assign _codeword[339] = message[309];
  assign _codeword[340] = message[310];
  assign _codeword[341] = message[311];
  assign _codeword[342] = message[312];
  assign _codeword[343] = message[313];
  assign _codeword[344] = message[314];
  assign _codeword[345] = message[315];
  assign _codeword[346] = message[316];
  assign _codeword[347] = message[317];
  assign _codeword[348] = message[318];
  assign _codeword[349] = message[319];
  assign _codeword[350] = message[320];
  assign _codeword[351] = message[321];
  assign _codeword[352] = message[322];
  assign _codeword[353] = message[323];
  assign _codeword[354] = message[324];
  assign _codeword[355] = message[325];
  assign _codeword[356] = message[326];
  assign _codeword[357] = message[327];
  assign _codeword[358] = message[328];
  assign _codeword[359] = message[329];
  assign _codeword[360] = message[330];
  assign _codeword[361] = message[331];
  assign _codeword[362] = message[332];
  assign _codeword[363] = message[333];
  assign _codeword[364] = message[334];
  assign _codeword[365] = message[335];
  assign _codeword[366] = message[336];
  assign _codeword[367] = message[337];
  assign _codeword[368] = message[338];
  assign _codeword[369] = message[339];
  assign _codeword[370] = message[340];
  assign _codeword[371] = message[341];
  assign _codeword[372] = message[342];
  assign _codeword[373] = message[343];
  assign _codeword[374] = message[344];
  assign _codeword[375] = message[345];
  assign _codeword[376] = message[346];
  assign _codeword[377] = message[347];
  assign _codeword[378] = message[348];
  assign _codeword[379] = message[349];
  assign _codeword[380] = message[350];
  assign _codeword[381] = message[351];
  assign _codeword[382] = message[352];
  assign _codeword[383] = message[353];
  assign _codeword[384] = message[354];
  assign _codeword[385] = message[355];
  assign _codeword[386] = message[356];
  assign _codeword[387] = message[357];
  assign _codeword[388] = message[358];
  assign _codeword[389] = message[359];
  assign _codeword[390] = message[360];
  assign _codeword[391] = message[361];
  assign _codeword[392] = message[362];
  assign _codeword[393] = message[363];
  assign _codeword[394] = message[364];
  assign _codeword[395] = message[365];
  assign _codeword[396] = message[366];
  assign _codeword[397] = message[367];
  assign _codeword[398] = message[368];
  assign _codeword[399] = message[369];
  assign _codeword[400] = message[370];
  assign _codeword[401] = message[371];
  assign _codeword[402] = message[372];
  assign _codeword[403] = message[373];
  assign _codeword[404] = message[374];
  assign _codeword[405] = message[375];
  assign _codeword[406] = message[376];
  assign _codeword[407] = message[377];
  assign _codeword[408] = message[378];
  assign _codeword[409] = message[379];
  assign _codeword[410] = message[380];
  assign _codeword[411] = message[381];
  assign _codeword[412] = message[382];
  assign _codeword[413] = message[383];
  assign _codeword[414] = message[384];
  assign _codeword[415] = message[385];
  assign _codeword[416] = message[386];
  assign _codeword[417] = message[387];
  assign _codeword[418] = message[388];
  assign _codeword[419] = message[389];
  assign _codeword[420] = message[390];
  assign _codeword[421] = message[391];
  assign _codeword[422] = message[392];
  assign _codeword[423] = message[393];
  assign _codeword[424] = message[394];
  assign _codeword[425] = message[395];
  assign _codeword[426] = message[396];
  assign _codeword[427] = message[397];
  assign _codeword[428] = message[398];
  assign _codeword[429] = message[399];
  assign _codeword[430] = message[400];
  assign _codeword[431] = message[401];
  assign _codeword[432] = message[402];
  assign _codeword[433] = message[403];
  assign _codeword[434] = message[404];
  assign _codeword[435] = message[405];
  assign _codeword[436] = message[406];
  assign _codeword[437] = message[407];
  assign _codeword[438] = message[408];
  assign _codeword[439] = message[409];
  assign _codeword[440] = message[410];
  assign _codeword[441] = message[411];
  assign _codeword[442] = message[412];
  assign _codeword[443] = message[413];
  assign _codeword[444] = message[414];
  assign _codeword[445] = message[415];
  assign _codeword[446] = message[416];
  assign _codeword[447] = message[417];
  assign _codeword[448] = message[418];
  assign _codeword[449] = message[419];
  assign _codeword[450] = message[420];
  assign _codeword[451] = message[421];
  assign _codeword[452] = message[422];
  assign _codeword[453] = message[423];
  assign _codeword[454] = message[424];
  assign _codeword[455] = message[425];
  assign _codeword[456] = message[426];
  assign _codeword[457] = message[427];
  assign _codeword[458] = message[428];
  assign _codeword[459] = message[429];
  assign _codeword[460] = message[430];
  assign _codeword[461] = message[431];
  assign _codeword[462] = message[432];
  assign _codeword[463] = message[433];
  assign _codeword[464] = message[434];
  assign _codeword[465] = message[435];
  assign _codeword[466] = message[436];
  assign _codeword[467] = message[437];
  assign _codeword[468] = message[438];
  assign _codeword[469] = message[439];
  assign _codeword[470] = message[440];
  assign _codeword[471] = message[441];
  assign _codeword[472] = message[442];
  assign _codeword[473] = message[443];
  assign _codeword[474] = message[444];
  assign _codeword[475] = message[445];
  assign _codeword[476] = message[446];
  assign _codeword[477] = message[447];
  assign _codeword[478] = message[448];
  assign _codeword[479] = message[449];
  assign _codeword[480] = message[450];
  assign _codeword[481] = message[451];
  assign _codeword[482] = message[452];
  assign _codeword[483] = message[453];
  assign _codeword[484] = message[454];
  assign _codeword[485] = message[455];
  assign _codeword[486] = message[456];
  assign _codeword[487] = message[457];
  assign _codeword[488] = message[458];
  assign _codeword[489] = message[459];
  assign _codeword[490] = message[460];
  assign _codeword[491] = message[461];
  assign _codeword[492] = message[462];
  assign _codeword[493] = message[463];
  assign _codeword[494] = message[464];
  assign _codeword[495] = message[465];
  assign _codeword[496] = message[466];
  assign _codeword[497] = message[467];
  assign _codeword[498] = message[468];
  assign _codeword[499] = message[469];
  assign _codeword[500] = message[470];
  assign _codeword[501] = message[471];
  assign _codeword[502] = message[472];
  assign _codeword[503] = message[473];
  assign _codeword[504] = message[474];
  assign _codeword[505] = message[475];
  assign _codeword[506] = message[476];
  assign _codeword[507] = message[477];
  assign _codeword[508] = message[478];
  assign _codeword[509] = message[479];
  assign _codeword[510] = message[480];
  assign _codeword[511] = message[481];
  assign _codeword[512] = message[482];
  assign _codeword[513] = message[483];
  assign _codeword[514] = message[484];
  assign _codeword[515] = message[485];
  assign _codeword[516] = message[486];
  assign _codeword[517] = message[487];
  assign _codeword[518] = message[488];
  assign _codeword[519] = message[489];
  assign _codeword[520] = message[490];
  assign _codeword[521] = message[491];
  assign _codeword[522] = message[492];
  assign _codeword[523] = message[493];
  assign _codeword[524] = message[494];
  assign _codeword[525] = message[495];
  assign _codeword[526] = message[496];
  assign _codeword[527] = message[497];
  assign _codeword[528] = message[498];
  assign _codeword[529] = message[499];
  assign _codeword[530] = message[500];
  assign _codeword[531] = message[501];
  assign _codeword[532] = message[502];
  assign _codeword[533] = message[503];
  assign _codeword[534] = message[504];
  assign _codeword[535] = message[505];
  assign _codeword[536] = message[506];
  assign _codeword[537] = message[507];
  assign _codeword[538] = message[508];
  assign _codeword[539] = message[509];
  assign _codeword[540] = message[510];
  assign _codeword[541] = message[511];

endmodule
