module GFDIV(a, b, c);
  input [7:0] a;
  input [7:0] b;
  output [7:0] c;

  /*
    GF(2^8)
    primitive polynomial : x^8 + x6 + x^4 + x^3 + x^2 + x + 1
    a = a^n
    b = a^m
    c = a/b = a^(n-m)
  */
  
  reg [7:0] binv;
  wire [7:0] imm;
  always_comb
      case (b)
        8'b0000_0000:  binv = 8'b0000_0000; // b=a^-inf => b=0 => a/0 = 0
        8'b0000_0001:  binv = 8'b0000_0001; // b=a^0 => a/(a^0) => a x (a^0)
        8'b0000_0010:  binv = 8'b1010_1111; // b=a^1 => a/(a^1) => a x (a^254)~~~~~
        8'b0000_0100:  binv = 8'b1111_1000; // b=a^2 
        8'b0000_1000:  binv = 8'b0111_1100; // b=a^3
        8'b0001_0000:  binv = 8'b0011_1110; // b=a^4 
        8'b0010_0000:  binv = 8'b0001_1111; // b=a^5 
        8'b0100_0000:  binv = 8'b1010_0000; // b=a^6 
        8'b1000_0000:  binv = 8'b0101_0000;//  b=a^7
        8'b0101_1111:  binv = 8'b0010_1000;//  b=a^8
        8'b1011_1110:  binv = 8'b0001_0100; // b=a^9
        8'b0010_0011:  binv = 8'b0000_1010; // b=a^10
        8'b0100_0110:  binv = 8'b0000_0101; // b=a^11
        8'b1000_1100:  binv = 8'b1010_1101; // b=a^12
        8'b0100_0111:  binv = 8'b1111_1001; // b=a^13
        8'b1000_1110:  binv = 8'b1101_0011; // b=a^14
        8'b0100_0011:  binv = 8'b1100_0110; // b=a^15
        8'b1000_0110:  binv = 8'b0110_0011; // b=a^16
        8'b0101_0011:  binv = 8'b1001_1110; // b=a^17
        8'b1010_0110:  binv = 8'b0100_1111; // b=a^18
        8'b0001_0011:  binv = 8'b1000_1000; // b=a^19
        8'b0010_0110:  binv = 8'b0100_0100; // b=a^20
        8'b0100_1100:  binv = 8'b0010_0010; // b=a^21
        8'b1001_1000:  binv = 8'b0001_0001; // b=a^22
        8'b0110_1111:  binv = 8'b1010_0111; // b=a^23
        8'b1101_1110:  binv = 8'b1111_1100; // b=a^24
        8'b1110_0011:  binv = 8'b0111_1110; // b=a^25
        8'b1001_1001:  binv = 8'b0011_1111; // b=a^26
        8'b0110_1101:  binv = 8'b1011_0000; // b=a^27
        8'b1101_1010:  binv = 8'b0101_1000; // b=a^28
        8'b1110_1011:  binv = 8'b0010_1100; // b=a^29
        8'b1000_1001:  binv = 8'b0001_0110; // b=a^30
        8'b0100_1101:  binv = 8'b0000_1011; // b=a^31
        8'b1001_1010:  binv = 8'b1010_1010; // b=a^32
        8'b0110_1011:  binv = 8'b0101_0101; // b=a^33
        8'b1101_0110:  binv = 8'b1000_0101; // b=a^34
        8'b1111_0011:  binv = 8'b1110_1101; // b=a^35
        8'b1011_1001:  binv = 8'b1101_1001; // b=a^36
        8'b0010_1101:  binv = 8'b1100_0011; // b=a^37
        8'b0101_1010:  binv = 8'b1100_1110; // b=a^38
        8'b1011_0100:  binv = 8'b0110_0111; // b=a^39
        8'b0011_0111:  binv = 8'b1001_1100; // b=a^40
        8'b0110_1110:  binv = 8'b0100_1110; // b=a^41
        8'b1101_1100:  binv = 8'b0010_0111; // b=a^42
        8'b1110_0111:  binv = 8'b1011_1100; // b=a^43
        8'b1001_0001:  binv = 8'b0101_1110; // b=a^44
        8'b0111_1101:  binv = 8'b0010_1111; // b=a^45
        8'b1111_1010:  binv = 8'b1011_1000; // b=a^46
        8'b1010_1011:  binv = 8'b0101_1100; // b=a^47
        8'b0000_1001:  binv = 8'b0010_1110; // b=a^48
        8'b0001_0010:  binv = 8'b0001_0111; // b=a^49
        8'b0010_0100:  binv = 8'b1010_0100; // b=a^50
        8'b0100_1000:  binv = 8'b0101_0010; // b=a^51
        8'b1001_0000:  binv = 8'b0010_1001; // b=a^52
        8'b0111_1111:  binv = 8'b1011_1011; // b=a^53
        8'b1111_1110:  binv = 8'b1111_0010; // b=a^54
        8'b1010_0011:  binv = 8'b0111_1001; // b=a^55
        8'b0001_1001:  binv = 8'b1001_0011; // b=a^56
        8'b0011_0010:  binv = 8'b1110_0110; // b=a^57
        8'b0110_0100:  binv = 8'b0111_0011; // b=a^58
        8'b1100_1000:  binv = 8'b1001_0110; // b=a^59
        8'b1100_1111:  binv = 8'b0100_1011; // b=a^60
        8'b1100_0001:  binv = 8'b1000_1010; // b=a^61
        8'b1101_1101:  binv = 8'b0100_0101; // b=a^62
        8'b1110_0101:  binv = 8'b1000_1101; // b=a^63
        8'b1001_0101:  binv = 8'b1110_1001; // b=a^64
        8'b0111_0101:  binv = 8'b1101_1011; // b=a^65
        8'b1110_1010:  binv = 8'b1100_0010; // b=a^66
        8'b1000_1011:  binv = 8'b0110_0001; // b=a^67
        8'b0100_1001:  binv = 8'b1001_1111; // b=a^68
        8'b1001_0010:  binv = 8'b1110_0000; // b=a^69
        8'b0111_1011:  binv = 8'b0111_0000; // b=a^70
        8'b1111_0110:  binv = 8'b0011_1000; // b=a^71
        8'b1011_0011:  binv = 8'b0001_1100; // b=a^72
        8'b0011_1001:  binv = 8'b0000_1110; // b=a^73
        8'b0111_0010:  binv = 8'b0000_0111; // b=a^74
        8'b1110_0100:  binv = 8'b1010_1100; // b=a^75
        8'b1001_0111:  binv = 8'b0101_0110; // b=a^76
        8'b0111_0001:  binv = 8'b0010_1011; // b=a^77
        8'b1110_0010:  binv = 8'b1011_1010; // b=a^78
        8'b1001_1011:  binv = 8'b0101_1101; // b=a^79
        8'b0110_1001:  binv = 8'b1000_0001; // b=a^80
        8'b1101_0010:  binv = 8'b1110_1111; // b=a^81
        8'b1111_1011:  binv = 8'b1101_1000; // b=a^82
        8'b1010_1001:  binv = 8'b0110_1100; // b=a^83
        8'b0000_1101:  binv = 8'b0011_0110; // b=a^84
        8'b0001_1010:  binv = 8'b0001_1011; // b=a^85
        8'b0011_0100:  binv = 8'b1010_0010; // b=a^86
        8'b0110_1000:  binv = 8'b0101_0001; // b=a^87
        8'b1101_0000:  binv = 8'b1000_0111; // b=a^88
        8'b1111_1111:  binv = 8'b1110_1100; // b=a^89
        8'b1010_0001:  binv = 8'b0111_0110; // b=a^90
        8'b0001_1101:  binv = 8'b0011_1011; // b=a^91
        8'b0011_1010:  binv = 8'b1011_0010; // b=a^92
        8'b0111_0100:  binv = 8'b0101_1001; // b=a^93
        8'b1110_1000:  binv = 8'b1000_0011; // b=a^94
        8'b1000_1111:  binv = 8'b1110_1110; // b=a^95
        8'b0100_0001:  binv = 8'b0111_0111; // b=a^96
        8'b1000_0010:  binv = 8'b1001_0100; // b=a^97
        8'b0101_1011:  binv = 8'b0100_1010; // b=a^98
        8'b1011_0110:  binv = 8'b0010_0101; // b=a^99
        8'b0011_0011:  binv = 8'b1011_1101; // b=a^100
        8'b0110_0110:  binv = 8'b1111_0001; // b=a^101
        8'b1100_1100:  binv = 8'b1101_0111; // b=a^102
        8'b1100_0111:  binv = 8'b1100_0100; // b=a^103
        8'b1101_0001:  binv = 8'b0110_0010; // b=a^104
        8'b1111_1101:  binv = 8'b0011_0001; // b=a^105
        8'b1010_0101:  binv = 8'b1011_0111; // b=a^106
        8'b0001_0101:  binv = 8'b1111_0100; // b=a^107
        8'b0010_1010:  binv = 8'b0111_1010; // b=a^108
        8'b0101_0100:  binv = 8'b0011_1101; // b=a^109
        8'b1010_1000:  binv = 8'b1011_0001; // b=a^110
        8'b0000_1111:  binv = 8'b1111_0111; // b=a^111
        8'b0001_1110:  binv = 8'b1101_0100; // b=a^112
        8'b0011_1100:  binv = 8'b0110_1010; // b=a^113
        8'b0111_1000:  binv = 8'b0011_0101; // b=a^114
        8'b1111_0000:  binv = 8'b1011_0101; // b=a^115
        8'b1011_1111:  binv = 8'b1111_0101; // b=a^116
        8'b0010_0001:  binv = 8'b1101_0101; // b=a^117
        8'b0100_0010:  binv = 8'b1100_0101; // b=a^118
        8'b1000_0100:  binv = 8'b1100_1101; // b=a^119
        8'b0101_0111:  binv = 8'b1100_1001; // b=a^120
        8'b1010_1110:  binv = 8'b1100_1011; // b=a^121
        8'b0000_0011:  binv = 8'b1100_1010; // b=a^122
        8'b0000_0110:  binv = 8'b0110_0101; // b=a^123
        8'b0000_1100:  binv = 8'b1001_1101; // b=a^124
        8'b0001_1000:  binv = 8'b1110_0001; // b=a^125
        8'b0011_0000:  binv = 8'b1101_1111; // b=a^126
        8'b0110_0000:  binv = 8'b1100_0000; // b=a^127
        8'b1100_0000:  binv = 8'b0110_0000; // b=a^128
        8'b1101_1111:  binv = 8'b0011_0000; // b=a^129
        8'b1110_0001:  binv = 8'b0001_1000; // b=a^130
        8'b1001_1101:  binv = 8'b0000_1100; // b=a^131
        8'b0110_0101:  binv = 8'b0000_0110; // b=a^132
        8'b1100_1010:  binv = 8'b0000_0011; // b=a^133
        8'b1100_1011:  binv = 8'b1010_1110; // b=a^134
        8'b1100_1001:  binv = 8'b0101_0111; // b=a^135
        8'b1100_1101:  binv = 8'b1000_0100; // b=a^136
        8'b1100_0101:  binv = 8'b0100_0010; // b=a^137
        8'b1101_0101:  binv = 8'b0010_0001; // b=a^138
        8'b1111_0101:  binv = 8'b1011_1111; // b=a^139
        8'b1011_0101:  binv = 8'b1111_0000; // b=a^140
        8'b0011_0101:  binv = 8'b0111_1000; // b=a^141
        8'b0110_1010:  binv = 8'b0011_1100; // b=a^142
        8'b1101_0100:  binv = 8'b0001_1110; // b=a^143
        8'b1111_0111:  binv = 8'b0000_1111; // b=a^144
        8'b1011_0001:  binv = 8'b1010_1000; // b=a^145
        8'b0011_1101:  binv = 8'b0101_0100; // b=a^146
        8'b0111_1010:  binv = 8'b0010_1010; // b=a^147
        8'b1111_0100:  binv = 8'b0001_0101; // b=a^148
        8'b1011_0111:  binv = 8'b1010_0101; // b=a^149
        8'b0011_0001:  binv = 8'b1111_1101; // b=a^150
        8'b0110_0010:  binv = 8'b1101_0001; // b=a^151
        8'b1100_0100:  binv = 8'b1100_0111; // b=a^152
        8'b1101_0111:  binv = 8'b1100_1100; // b=a^153
        8'b1111_0001:  binv = 8'b0110_0110; // b=a^154
        8'b1011_1101:  binv = 8'b0011_0011; // b=a^155
        8'b0010_0101:  binv = 8'b1011_0110; // b=a^156
        8'b0100_1010:  binv = 8'b0101_1011; // b=a^157
        8'b1001_0100:  binv = 8'b1000_0010; // b=a^158
        8'b0111_0111:  binv = 8'b0100_0001; // b=a^159
        8'b1110_1110:  binv = 8'b1000_1111; // b=a^160
        8'b1000_0011:  binv = 8'b1110_1000; // b=a^161
        8'b0101_1001:  binv = 8'b0111_0100; // b=a^162
        8'b1011_0010:  binv = 8'b0011_1010; // b=a^163
        8'b0011_1011:  binv = 8'b0001_1101; // b=a^164
        8'b0111_0110:  binv = 8'b1010_0001; // b=a^165
        8'b1110_1100:  binv = 8'b1111_1111; // b=a^166 
        8'b1000_0111:  binv = 8'b1101_0000; // b=a^167
        8'b0101_0001:  binv = 8'b0110_1000; // b=a^168
        8'b1010_0010:  binv = 8'b0011_0100; // b=a^169
        8'b0001_1011:  binv = 8'b0001_1010; // b=a^170
        8'b0011_0110:  binv = 8'b0000_1101; // b=a^171
        8'b0110_1100:  binv = 8'b1010_1001; // b=a^172
        8'b1101_1000:  binv = 8'b1111_1011; // b=a^173
        8'b1110_1111:  binv = 8'b1101_0010; // b=a^174
        8'b1000_0001:  binv = 8'b0110_1001; // b=a^175
        8'b0101_1101:  binv = 8'b1001_1011; // b=a^176
        8'b1011_1010:  binv = 8'b1110_0010; // b=a^177
        8'b0010_1011:  binv = 8'b0111_0001; // b=a^178
        8'b0101_0110:  binv = 8'b1001_0111; // b=a^179
        8'b1010_1100:  binv = 8'b1110_0100; // b=a^180
        8'b0000_0111:  binv = 8'b0111_0010; // b=a^181
        8'b0000_1110:  binv = 8'b0011_1001; // b=a^182
        8'b0001_1100:  binv = 8'b1011_0011; // b=a^183
        8'b0011_1000:  binv = 8'b1111_0110; // b=a^184
        8'b0111_0000:  binv = 8'b0111_1011; // b=a^185
        8'b1110_0000:  binv = 8'b1001_0010; // b=a^186
        8'b1001_1111:  binv = 8'b0100_1001; // b=a^187
        8'b0110_0001:  binv = 8'b1000_1011; // b=a^188
        8'b1100_0010:  binv = 8'b1110_1010; // b=a^189
        8'b1101_1011:  binv = 8'b0111_0101; // b=a^190
        8'b1110_1001:  binv = 8'b1001_0101; // b=a^191
        8'b1000_1101:  binv = 8'b1110_0101; // b=a^192
        8'b0100_0101:  binv = 8'b1101_1101; // b=a^193
        8'b1000_1010:  binv = 8'b1100_0001; // b=a^194
        8'b0100_1011:  binv = 8'b1100_1111; // b=a^195
        8'b1001_0110:  binv = 8'b1100_1000; // b=a^196
        8'b0111_0011:  binv = 8'b0110_0100; // b=a^197
        8'b1110_0110:  binv = 8'b0011_0010; // b=a^198
        8'b1001_0011:  binv = 8'b0001_1001; // b=a^199
        8'b0111_1001:  binv = 8'b1010_0011; // b=a^200
        8'b1111_0010:  binv = 8'b1111_1110; // b=a^201
        8'b1011_1011:  binv = 8'b0111_1111; // b=a^202
        8'b0010_1001:  binv = 8'b1001_0000; // b=a^203
        8'b0101_0010:  binv = 8'b0100_1000; // b=a^204
        8'b1010_0100:  binv = 8'b0010_0100; // b=a^205
        8'b0001_0111:  binv = 8'b0001_0010; // b=a^206
        8'b0010_1110:  binv = 8'b0000_1001; // b=a^207
        8'b0101_1100:  binv = 8'b1010_1011; // b=a^208
        8'b1011_1000:  binv = 8'b1111_1010; // b=a^209
        8'b0010_1111:  binv = 8'b0111_1101; // b=a^210
        8'b0101_1110:  binv = 8'b1001_0001; // b=a^211
        8'b1011_1100:  binv = 8'b1110_0111; // b=a^212
        8'b0010_0111:  binv = 8'b1101_1100; // b=a^213
        8'b0100_1110:  binv = 8'b0110_1110; // b=a^214
        8'b1001_1100:  binv = 8'b0011_0111; // b=a^215
        8'b0110_0111:  binv = 8'b1011_0100; // b=a^216
        8'b1100_1110:  binv = 8'b0101_1010; // b=a^217
        8'b1100_0011:  binv = 8'b0010_1101; // b=a^218
        8'b1101_1001:  binv = 8'b1011_1001; // b=a^219
        8'b1110_1101:  binv = 8'b1111_0011; // b=a^220
        8'b1000_0101:  binv = 8'b1101_0110; // b=a^221
        8'b0101_0101:  binv = 8'b0110_1011; // b=a^222
        8'b1010_1010:  binv = 8'b1001_1010; // b=a^223
        8'b0000_1011:  binv = 8'b0100_1101; // b=a^224
        8'b0001_0110:  binv = 8'b1000_1001; // b=a^225
        8'b0010_1100:  binv = 8'b1110_1011; // b=a^226
        8'b0101_1000:  binv = 8'b1101_1010; // b=a^227
        8'b1011_0000:  binv = 8'b0110_1101; // b=a^228
        8'b0011_1111:  binv = 8'b1001_1001; // b=a^229
        8'b0111_1110:  binv = 8'b1110_0011; // b=a^230
        8'b1111_1100:  binv = 8'b1101_1110; // b=a^231
        8'b1010_0111:  binv = 8'b0110_1111; // b=a^232
        8'b0001_0001:  binv = 8'b1001_1000; // b=a^233
        8'b0010_0010:  binv = 8'b0100_1100; // b=a^234
        8'b0100_0100:  binv = 8'b0010_0110; // b=a^235
        8'b1000_1000:  binv = 8'b0001_0011; // b=a^236
        8'b0100_1111:  binv = 8'b1010_0110; // b=a^237
        8'b1001_1110:  binv = 8'b0101_0011; // b=a^238
        8'b0110_0011:  binv = 8'b1000_0110; // b=a^239
        8'b1100_0110:  binv = 8'b0100_0011; // b=a^240
        8'b1101_0011:  binv = 8'b1000_1110; // b=a^241
        8'b1111_1001:  binv = 8'b0100_0111; // b=a^242
        8'b1010_1101:  binv = 8'b1000_1100; // b=a^243
        8'b0000_0101:  binv = 8'b0100_0110; // b=a^244
        8'b0000_1010:  binv = 8'b0010_0011; // b=a^245
        8'b0001_0100:  binv = 8'b1011_1110; // b=a^246
        8'b0010_1000:  binv = 8'b0101_1111; // b=a^247
        8'b0101_0000:  binv = 8'b1000_0000; // b=a^248
        8'b1010_0000:  binv = 8'b0100_0000; // b=a^249
        8'b0001_1111:  binv = 8'b0010_0000; // b=a^250
        8'b0011_1110:  binv = 8'b0001_0000; // b=a^251
        8'b0111_1100:  binv = 8'b0000_1000; // b=a^252
        8'b1111_1000:  binv = 8'b0000_0100; // b=a^253
        8'b1010_1111:  binv = 8'b0000_0010; // b=a^254
      endcase
    GFMULT gfmult(a, binv, imm);
    assign c = imm;

endmodule

