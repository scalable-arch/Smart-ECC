module encoder_tb;
  reg [511:0] message;
  wire [541:0] codeword;
  integer failures;

  bch_encoder encoder(message, codeword);

  initial
  begin
    failures = 0;

    message <= 512'b11011001110110100111101111101010000110100011000111011000101010111110001010100010011110110100111010000101010111000101110001011100010100001110110100000000110001001000001110001000111010101001101100001111101101111100001000000100110000101100000100101101001110011001011100010101011110100110111111001000111001001011101111100100001100101100010000001101001101011111001001110001011000001001001011101011101000000010111000110111100110000001011111010110001101101010000101000100010101010001110111110100100110101101111000110111;
    #1;
    if (codeword != 542'b11011001110110100111101111101010000110100011000111011000101010111110001010100010011110110100111010000101010111000101110001011100010100001110110100000000110001001000001110001000111010101001101100001111101101111100001000000100110000101100000100101101001110011001011100010101011110100110111111001000111001001011101111100100001100101100010000001101001101011111001001110001011000001001001011101011101000000010111000110111100110000001011111010110001101101010000101000100010101010001110111110100100110101101111000110111100100010111011011110010010001)
      failures = failures+1;

    message <= 512'b11110000000111110010111001110010010010101100000010101011001101011011111000111010001000001111111101111010011111010111111111001010110100000000010110100011001100100001101110111111000010000101110000101011110001100001000110101110100010000010000010000011100111010010011111101100101100101110001110100101111011100011100010010100100010000101101101010010100010010011000001110100000000001110001110011000010101000110101110000011000000111001111010001001111011101101010000011101110010011110010111111001101011000001011101010001;
    #1;
    if (codeword != 542'b11110000000111110010111001110010010010101100000010101011001101011011111000111010001000001111111101111010011111010111111111001010110100000000010110100011001100100001101110111111000010000101110000101011110001100001000110101110100010000010000010000011100111010010011111101100101100101110001110100101111011100011100010010100100010000101101101010010100010010011000001110100000000001110001110011000010101000110101110000011000000111001111010001001111011101101010000011101110010011110010111111001101011000001011101010001101000111010001110011011111111)
      failures = failures+1;

    message <= 512'b00101010111101110000110101101011111100000110011111010011011111101101010000011101110011001010011100000100110000111000101101001111010111011011101010011011100100111100001101010101101001010111011001100000000010100011111000011110110111100101110000111001011011111111001101110111101001110101110001111101001110110001011001111001110100010000110011110100000001001111111000010010111100111111000111101101101100011011110010001010110101100000111101010101111100111011011011011110011000001000000000000101000000000011100010000010;
    #1;
    if (codeword != 542'b00101010111101110000110101101011111100000110011111010011011111101101010000011101110011001010011100000100110000111000101101001111010111011011101010011011100100111100001101010101101001010111011001100000000010100011111000011110110111100101110000111001011011111111001101110111101001110101110001111101001110110001011001111001110100010000110011110100000001001111111000010010111100111111000111101101101100011011110010001010110101100000111101010101111100111011011011011110011000001000000000000101000000000011100010000010001111010010100001001100011011)
      failures = failures+1;

    message <= 512'b11011110100110011110101011000001010000111100000111001111110100001010010110011100111110100101100010000000010110010010111101011100011110110100101111110010001110011100111010100011000110001100100101110110100011010110101001100101110011111010001111111000111101101000010000010001011011011001110111100000011000000101000001011100011001101101001101110001001100010010110011110100011110101110011111110100100100000100001011110010111010001111010111110010000111011110101110100110110000010101011000000111010110111110001100111011;
    #1;
    if (codeword != 542'b11011110100110011110101011000001010000111100000111001111110100001010010110011100111110100101100010000000010110010010111101011100011110110100101111110010001110011100111010100011000110001100100101110110100011010110101001100101110011111010001111111000111101101000010000010001011011011001110111100000011000000101000001011100011001101101001101110001001100010010110011110100011110101110011111110100100100000100001011110010111010001111010111110010000111011110101110100110110000010101011000000111010110111110001100111011100001110010100101001111000000)
      failures = failures+1;

    message <= 512'b00011011001111001110111011011010100100001100101111011111011001011110011111101101101000001000101110110001011100100001111000110001100010101111101000101111011101110001110111001110011000111101100001111010000101110111010010001001011101010101100011011000100001111101000110010110011101011001001011111010111001111000000100000100001101011101001101101000100101111001101111110010101001011001000001000101000110111110000100010011000101011010110011001011011100111101111010111111000000011001001101100100011001010000001011110011;
    #1;
    if (codeword != 542'b00011011001111001110111011011010100100001100101111011111011001011110011111101101101000001000101110110001011100100001111000110001100010101111101000101111011101110001110111001110011000111101100001111010000101110111010010001001011101010101100011011000100001111101000110010110011101011001001011111010111001111000000100000100001101011101001101101000100101111001101111110010101001011001000001000101000110111110000100010011000101011010110011001011011100111101111010111111000000011001001101100100011001010000001011110011001011001110101001010011111111)
      failures = failures+1;

    message <= 512'b10010111100001100100101001111001011010110110111100101110010101011100110110100110100000000010100001011111111001101000000011100111111111100100010110001100111101101100010010011010010011100010010111111000110010000000100110000101111111000101111100100011101101011001010011110111101110010011000111100001111110100110011000000100110010111001101011101010010111000010110111100100111101111011101010010110001011110011001010011101011101110010011110010101001100110010000101001001001110000110101011100001011110011010101000100110;
    #1;
    if (codeword != 542'b10010111100001100100101001111001011010110110111100101110010101011100110110100110100000000010100001011111111001101000000011100111111111100100010110001100111101101100010010011010010011100010010111111000110010000000100110000101111111000101111100100011101101011001010011110111101110010011000111100001111110100110011000000100110010111001101011101010010111000010110111100100111101111011101010010110001011110011001010011101011101110010011110010101001100110010000101001001001110000110101011100001011110011010101000100110011101100110111011001111101101)
      failures = failures+1;

    message <= 512'b01101000000001100100101001101101110000100010100010011011001100111011100011011100110010110001110110011100010001011110111111000001000110011111101011100000001111010011011000110110011000001000101000101001011111001011110011111110101010011111111110101001110110110100011111110100001100100110001110101100010001110010100011100001111010111001111111010010101001000001111011101000110001011001100010100011011110001010110101000001100110111100100011111011000000000111111101010000110111011101011101100100111000111001011101010010;
    #1;
    if (codeword != 542'b01101000000001100100101001101101110000100010100010011011001100111011100011011100110010110001110110011100010001011110111111000001000110011111101011100000001111010011011000110110011000001000101000101001011111001011110011111110101010011111111110101001110110110100011111110100001100100110001110101100010001110010100011100001111010111001111111010010101001000001111011101000110001011001100010100011011110001010110101000001100110111100100011111011000000000111111101010000110111011101011101100100111000111001011101010010000100011010011000000111100111)
      failures = failures+1;

    message <= 512'b00100100110110111111000010100111001011011100001101100100110100110110110100010000111100111000010010011101011100010010111001011111111000101101111101100101001010011111110010011010000001100000000111110111010110100000111111111101011100011001110010001010111101000100010011100111000111000011111110101001011010110000010101011101110010001101111110101101000110110011100001011011010111001001110011000110110010110001001101000001011111011011101100110001010101011001000001011001011101000111101100011011100011000011011101010110;
    #1;
    if (codeword != 542'b00100100110110111111000010100111001011011100001101100100110100110110110100010000111100111000010010011101011100010010111001011111111000101101111101100101001010011111110010011010000001100000000111110111010110100000111111111101011100011001110010001010111101000100010011100111000111000011111110101001011010110000010101011101110010001101111110101101000110110011100001011011010111001001110011000110110010110001001101000001011111011011101100110001010101011001000001011001011101000111101100011011100011000011011101010110000100000000001000000100001001)
      failures = failures+1;

    message <= 512'b10001100011010011100000110111000010111001010110000110001111101001010010101100010001010010100111001100111001010010110000110001111101000001100000010001111110110100001100011001110110010011111000010001111110110011011000000010000001010010010111111110110101111101011101010111001111010110101000010000011000001001101001110010010100001100001011100100110001101101011001111110001101010111001000101001100010101000111111110011010000101010111111001000101110010000110001100111001000111000001111111100000110010000110110100011111;
    #1;
    if (codeword != 542'b10001100011010011100000110111000010111001010110000110001111101001010010101100010001010010100111001100111001010010110000110001111101000001100000010001111110110100001100011001110110010011111000010001111110110011011000000010000001010010010111111110110101111101011101010111001111010110101000010000011000001001101001110010010100001100001011100100110001101101011001111110001101010111001000101001100010101000111111110011010000101010111111001000101110010000110001100111001000111000001111111100000110010000110110100011111000101100011001010010100001110)
      failures = failures+1;

    message <= 512'b00001010010101010100010011011010011011000010111011000110011001111011011011011110101100100100011101011011100100101110101101100100011011000101001101011111011100000011011111010010001111110110010101011001001011011111100000111100010111010011010000010100100111101010011001001111111110100010011000011110101100010000010101001110100000000011011100110011101100010011001010111011101101010001001101101010010110010100010011100100110101001001001000000110011110100010110111001101010110001111011010001110000100100111111001111000;
    #1;
    if (codeword != 542'b00001010010101010100010011011010011011000010111011000110011001111011011011011110101100100100011101011011100100101110101101100100011011000101001101011111011100000011011111010010001111110110010101011001001011011111100000111100010111010011010000010100100111101010011001001111111110100010011000011110101100010000010101001110100000000011011100110011101100010011001010111011101101010001001101101010010110010100010011100100110101001001001000000110011110100010110111001101010110001111011010001110000100100111111001111000100011010000101011100100001101)
      failures = failures+1;

    message <= 512'b01011101001101010001111101010110100111000011011111001011010010000110111101111110000011110000000000101001111111001010001111111000110100111111001000111111010001110110011000101101111000000101100010100111001100010000000010100110001110110101110101110001101000111000010010111011101011010101110011001101110001010011100011111100110000010010000010111111010000010111000100011101001011000010101000001001000010110010001101001000101001011110001010011100011111011110101101011100110101100100001010000101001011000100110101110011;
    #1;
    if (codeword != 542'b01011101001101010001111101010110100111000011011111001011010010000110111101111110000011110000000000101001111111001010001111111000110100111111001000111111010001110110011000101101111000000101100010100111001100010000000010100110001110110101110101110001101000111000010010111011101011010101110011001101110001010011100011111100110000010010000010111111010000010111000100011101001011000010101000001001000010110010001101001000101001011110001010011100011111011110101101011100110101100100001010000101001011000100110101110011011100011001010111001110010101)
      failures = failures+1;

    message <= 512'b00000001110100110000000110101100010111000100110100111001101001010000111111000010101101001001011011011110101101100111001101110000010011011100000010010011010110000011010111010001000111100101100011010110011100110110000010110110101001111010001111100010100001111110000000100001001000100101101111100111010111011000110100001001101011001100011100100010011101110101100000101111011111100101010101001001011110001000000011000001101000111000010010001101101101001011110110000011010010000101100101101010101111100010011010000000;
    #1;
    if (codeword != 542'b00000001110100110000000110101100010111000100110100111001101001010000111111000010101101001001011011011110101101100111001101110000010011011100000010010011010110000011010111010001000111100101100011010110011100110110000010110110101001111010001111100010100001111110000000100001001000100101101111100111010111011000110100001001101011001100011100100010011101110101100000101111011111100101010101001001011110001000000011000001101000111000010010001101101101001011110110000011010010000101100101101010101111100010011010000000010001001110111111011000001101)
      failures = failures+1;

    message <= 512'b11011111011001001000010110101011001111010101111011101001111111110001100001111100011000111011011000101001111110100011111111010110111011100000010101111101011000111000000101100110111101100111110000110001010110000001011111110111101111011010011010000000011000010101111110100000000111011101011101110000001101110101101100000101011100000000010011000000011100000100100001101011001000011101100110101101001111000011000101011100110111110010010101100101101111101111110100001011110010001010000110100111011110010001111110011111;
    #1;
    if (codeword != 542'b11011111011001001000010110101011001111010101111011101001111111110001100001111100011000111011011000101001111110100011111111010110111011100000010101111101011000111000000101100110111101100111110000110001010110000001011111110111101111011010011010000000011000010101111110100000000111011101011101110000001101110101101100000101011100000000010011000000011100000100100001101011001000011101100110101101001111000011000101011100110111110010010101100101101111101111110100001011110010001010000110100111011110010001111110011111101100100000011111011000111000)
      failures = failures+1;

    message <= 512'b00101100111101011101100111110110010011101010110010111111001010110000110010101010011010111011000010110101010100011110100101011001000001110010011010110110000110101001110101101100011100111110111111000011010000001111001011010110011111111000111010101101001000111001000011000010100110111000000010110111000001000010001011010111000111011010110110010110111110000000011101101010101010010111100011011000110101111010010010100110001001110111101000001100000011100011100011000111100010001101110110001000010100001101010101000101;
    #1;
    if (codeword != 542'b00101100111101011101100111110110010011101010110010111111001010110000110010101010011010111011000010110101010100011110100101011001000001110010011010110110000110101001110101101100011100111110111111000011010000001111001011010110011111111000111010101101001000111001000011000010100110111000000010110111000001000010001011010111000111011010110110010110111110000000011101101010101010010111100011011000110101111010010010100110001001110111101000001100000011100011100011000111100010001101110110001000010100001101010101000101101100101010011001100110011110)
      failures = failures+1;

    message <= 512'b00100011001010011011111000001011101001101010111010110011110000001111100100101010110001101110101100010100111100101011001000100100001110010000101000111000001011010001110101110011000100100111001100000000010011000010011011110100000110100101110010101101110010011110001111100100100010001000001111101111000100101101100100101000010101010111001100011011000010011011101010000001110101001011100011111110111110000001011010110110101011010110100101100010101100101110111111100001000010000101101101010010000011110101010100001010;
    #1;
    if (codeword != 542'b00100011001010011011111000001011101001101010111010110011110000001111100100101010110001101110101100010100111100101011001000100100001110010000101000111000001011010001110101110011000100100111001100000000010011000010011011110100000110100101110010101101110010011110001111100100100010001000001111101111000100101101100100101000010101010111001100011011000010011011101010000001110101001011100011111110111110000001011010110110101011010110100101100010101100101110111111100001000010000101101101010010000011110101010100001010010100110011011000100111110001)
      failures = failures+1;

    message <= 512'b10011111101001001000110001000111000111110111000101100110011010000110000101110110110110011110001101000100101111110111010100101110101010100011010010101111001010110011110101011001001111110101100010011100011110000001100101101110110111000011000000010100101101110101101100011000111001110111101000001000010110001010100011110110100001001111000110111011111100010100011100011110110001100111110011010101100111111101011100011110001001111101101101010011111100110110110101101111000110101001000011111010010000101011101000000000;
    #1;
    if (codeword != 542'b10011111101001001000110001000111000111110111000101100110011010000110000101110110110110011110001101000100101111110111010100101110101010100011010010101111001010110011110101011001001111110101100010011100011110000001100101101110110111000011000000010100101101110101101100011000111001110111101000001000010110001010100011110110100001001111000110111011111100010100011100011110110001100111110011010101100111111101011100011110001001111101101101010011111100110110110101101111000110101001000011111010010000101011101000000000001010010111001101010010111000)
      failures = failures+1;

    message <= 512'b10101101011011010101001000011110010101110001010110000001100111110100111100010010011100011100010100111101100011101001100001010000000000010101111100001011100101110010111111101010011011110001100000010001111100011000100010000101010011101011100010110000001110101111011010011010001010111011001010111100100000101101001001110010111000100101001111000101011100101001010010011110110000101010111010011010000010101100100111101110111111000111000100010110000100110100111010011110100100101001000111001011101110000001100110010001;
    #1;
    if (codeword != 542'b10101101011011010101001000011110010101110001010110000001100111110100111100010010011100011100010100111101100011101001100001010000000000010101111100001011100101110010111111101010011011110001100000010001111100011000100010000101010011101011100010110000001110101111011010011010001010111011001010111100100000101101001001110010111000100101001111000101011100101001010010011110110000101010111010011010000010101100100111101110111111000111000100010110000100110100111010011110100100101001000111001011101110000001100110010001000101110010000000000111110110)
      failures = failures+1;

    message <= 512'b01000011000100110101011101011011001000110000011111000000010101100001100010100101011010111101000011010001110101100001000111000101111010001100000001000011100110100001010001010010001001000011111110010000110100011001111100100111110110110011100010000110111111001000110101110100110110100010001000000111110100100000011011001101001111110010100010010111011101001111010000001010111101000010110000010000001010011001000001110000100101111111000011000010101011010011110100100100100000100011111111111010100010010011111111000101;
    #1;
    if (codeword != 542'b01000011000100110101011101011011001000110000011111000000010101100001100010100101011010111101000011010001110101100001000111000101111010001100000001000011100110100001010001010010001001000011111110010000110100011001111100100111110110110011100010000110111111001000110101110100110110100010001000000111110100100000011011001101001111110010100010010111011101001111010000001010111101000010110000010000001010011001000001110000100101111111000011000010101011010011110100100100100000100011111111111010100010010011111111000101110100001000111111000010101001)
      failures = failures+1;

    message <= 512'b11010111011001010010010110011100000111001010110011010010011110110010000011101110001011010101101111000110110000000011101111101110110110001101101110011000001010110101111010111110101110110001110100110000000011011011010010111110111101011000111001101101000011011000110101011100011101100101010001000101101001111100101111010100001101101000110110100000011010110111100001001100001011100000011110001101111010110001101111101111000011010111100000010111010011011000011111100011111110110111111111010101001111111100101100111100;
    #1;
    if (codeword != 542'b11010111011001010010010110011100000111001010110011010010011110110010000011101110001011010101101111000110110000000011101111101110110110001101101110011000001010110101111010111110101110110001110100110000000011011011010010111110111101011000111001101101000011011000110101011100011101100101010001000101101001111100101111010100001101101000110110100000011010110111100001001100001011100000011110001101111010110001101111101111000011010111100000010111010011011000011111100011111110110111111111010101001111111100101100111100001111000101101100111000010010)
      failures = failures+1;

    message <= 512'b00011101011100101110011110110111011011100100010111001111100001000100000110001110001010100011011010011110110110010001011100111111111111101001000010001001001111110101001010011101000111100010000001110101010101100000001000000101011110101100010000110000000110011100101110101100011000100000100000001101000110000011111111010000000110100111100001010011110010110100011111101100101010010110000110110111001000010101001101110000000110100100000001010011010001000001111011000111011111111110110010110011111010110101111100011110;
    #1;
    if (codeword != 542'b00011101011100101110011110110111011011100100010111001111100001000100000110001110001010100011011010011110110110010001011100111111111111101001000010001001001111110101001010011101000111100010000001110101010101100000001000000101011110101100010000110000000110011100101110101100011000100000100000001101000110000011111111010000000110100111100001010011110010110100011111101100101010010110000110110111001000010101001101110000000110100100000001010011010001000001111011000111011111111110110010110011111010110101111100011110101001000101001111001011110001)
      failures = failures+1;

    $display("\n==============================");
    if (!failures)
      $display("\nAll encoding tests passed\n");
    else
      $display("Failed %d encoding test(s)", failures);
    $display("==============================\n");
  end
endmodule
