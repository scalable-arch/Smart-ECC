module bch_syndromes(received, syndrome1, syndrome2, syndrome3, syndrome4, syndrome5);
  input [541:0] received;
  output [9:0] syndrome1;
  output [9:0] syndrome2;
  output [9:0] syndrome3;
  output [9:0] syndrome4;
  output [9:0] syndrome5;

  assign syndrome1 = ({10{received[0]}} & 10'b0000000001) ^ 
  ({10{received[1]}} & 10'b0000000010) ^ ({10{received[2]}} & 10'b0000000100) ^ ({10{received[3]}} & 10'b0000001000) ^ ({10{received[4]}} & 10'b0000010000) ^ ({10{received[5]}} & 10'b0000100000) ^ ({10{received[6]}} & 10'b0001000000) ^ ({10{received[7]}} & 10'b0010000000) ^ ({10{received[8]}} & 10'b0100000000) ^ ({10{received[9]}} & 10'b1000000000) ^ ({10{received[10]}} & 10'b0000001001) ^ ({10{received[11]}} & 10'b0000010010) ^ ({10{received[12]}} & 10'b0000100100) ^ ({10{received[13]}} & 10'b0001001000) ^ ({10{received[14]}} & 10'b0010010000) ^ ({10{received[15]}} & 10'b0100100000) ^ ({10{received[16]}} & 10'b1001000000) ^ ({10{received[17]}} & 10'b0010001001) ^ ({10{received[18]}} & 10'b0100010010) ^ ({10{received[19]}} & 10'b1000100100) ^ ({10{received[20]}} & 10'b0001000001) ^ ({10{received[21]}} & 10'b0010000010) ^ ({10{received[22]}} & 10'b0100000100) ^ ({10{received[23]}} & 10'b1000001000) ^ ({10{received[24]}} & 10'b0000011001) ^ ({10{received[25]}} & 10'b0000110010) ^ ({10{received[26]}} & 10'b0001100100) ^ ({10{received[27]}} & 10'b0011001000) ^ ({10{received[28]}} & 10'b0110010000) ^ ({10{received[29]}} & 10'b1100100000) ^ ({10{received[30]}} & 10'b1001001001) ^ ({10{received[31]}} & 10'b0010011011) ^ ({10{received[32]}} & 10'b0100110110) ^ ({10{received[33]}} & 10'b1001101100) ^ ({10{received[34]}} & 10'b0011010001) ^ ({10{received[35]}} & 10'b0110100010) ^ ({10{received[36]}} & 10'b1101000100) ^ ({10{received[37]}} & 10'b1010000001) ^ ({10{received[38]}} & 10'b0100001011) ^ ({10{received[39]}} & 10'b1000010110) ^ ({10{received[40]}} & 10'b0000100101) ^ ({10{received[41]}} & 10'b0001001010) ^ ({10{received[42]}} & 10'b0010010100) ^ ({10{received[43]}} & 10'b0100101000) ^ ({10{received[44]}} & 10'b1001010000) ^ ({10{received[45]}} & 10'b0010101001) ^ ({10{received[46]}} & 10'b0101010010) ^ ({10{received[47]}} & 10'b1010100100) ^ ({10{received[48]}} & 10'b0101000001) ^ ({10{received[49]}} & 10'b1010000010) ^ ({10{received[50]}} & 10'b0100001101) ^ ({10{received[51]}} & 10'b1000011010) ^ ({10{received[52]}} & 10'b0000111101) ^ ({10{received[53]}} & 10'b0001111010) ^ ({10{received[54]}} & 10'b0011110100) ^ ({10{received[55]}} & 10'b0111101000) ^ ({10{received[56]}} & 10'b1111010000) ^ ({10{received[57]}} & 10'b1110101001) ^ ({10{received[58]}} & 10'b1101011011) ^ ({10{received[59]}} & 10'b1010111111) ^ ({10{received[60]}} & 10'b0101110111) ^ ({10{received[61]}} & 10'b1011101110) ^ ({10{received[62]}} & 10'b0111010101) ^ ({10{received[63]}} & 10'b1110101010) ^ ({10{received[64]}} & 10'b1101011101) ^ ({10{received[65]}} & 10'b1010110011) ^ ({10{received[66]}} & 10'b0101101111) ^ ({10{received[67]}} & 10'b1011011110) ^ ({10{received[68]}} & 10'b0110110101) ^ ({10{received[69]}} & 10'b1101101010) ^ ({10{received[70]}} & 10'b1011011101) ^ ({10{received[71]}} & 10'b0110110011) ^ ({10{received[72]}} & 10'b1101100110) ^ ({10{received[73]}} & 10'b1011000101) ^ ({10{received[74]}} & 10'b0110000011) ^ ({10{received[75]}} & 10'b1100000110) ^ ({10{received[76]}} & 10'b1000000101) ^ ({10{received[77]}} & 10'b0000000011) ^ ({10{received[78]}} & 10'b0000000110) ^ ({10{received[79]}} & 10'b0000001100) ^ ({10{received[80]}} & 10'b0000011000) ^ ({10{received[81]}} & 10'b0000110000) ^ ({10{received[82]}} & 10'b0001100000) ^ ({10{received[83]}} & 10'b0011000000) ^ ({10{received[84]}} & 10'b0110000000) ^ ({10{received[85]}} & 10'b1100000000) ^ ({10{received[86]}} & 10'b1000001001) ^ ({10{received[87]}} & 10'b0000011011) ^ ({10{received[88]}} & 10'b0000110110) ^ ({10{received[89]}} & 10'b0001101100) ^ ({10{received[90]}} & 10'b0011011000) ^ ({10{received[91]}} & 10'b0110110000) ^ ({10{received[92]}} & 10'b1101100000) ^ ({10{received[93]}} & 10'b1011001001) ^ ({10{received[94]}} & 10'b0110011011) ^ ({10{received[95]}} & 10'b1100110110) ^ ({10{received[96]}} & 10'b1001100101) ^ ({10{received[97]}} & 10'b0011000011) ^ ({10{received[98]}} & 10'b0110000110) ^ ({10{received[99]}} & 10'b1100001100) ^ ({10{received[100]}} & 10'b1000010001) ^ ({10{received[101]}} & 10'b0000101011) ^ ({10{received[102]}} & 10'b0001010110) ^ ({10{received[103]}} & 10'b0010101100) ^ ({10{received[104]}} & 10'b0101011000) ^ ({10{received[105]}} & 10'b1010110000) ^ ({10{received[106]}} & 10'b0101101001) ^ ({10{received[107]}} & 10'b1011010010) ^ ({10{received[108]}} & 10'b0110101101) ^ ({10{received[109]}} & 10'b1101011010) ^ ({10{received[110]}} & 10'b1010111101) ^ ({10{received[111]}} & 10'b0101110011) ^ ({10{received[112]}} & 10'b1011100110) ^ ({10{received[113]}} & 10'b0111000101) ^ ({10{received[114]}} & 10'b1110001010) ^ ({10{received[115]}} & 10'b1100011101) ^ ({10{received[116]}} & 10'b1000110011) ^ ({10{received[117]}} & 10'b0001101111) ^ ({10{received[118]}} & 10'b0011011110) ^ ({10{received[119]}} & 10'b0110111100) ^ ({10{received[120]}} & 10'b1101111000) ^ ({10{received[121]}} & 10'b1011111001) ^ ({10{received[122]}} & 10'b0111111011) ^ ({10{received[123]}} & 10'b1111110110) ^ ({10{received[124]}} & 10'b1111100101) ^ ({10{received[125]}} & 10'b1111000011) ^ ({10{received[126]}} & 10'b1110001111) ^ ({10{received[127]}} & 10'b1100010111) ^ ({10{received[128]}} & 10'b1000100111) ^ ({10{received[129]}} & 10'b0001000111) ^ ({10{received[130]}} & 10'b0010001110) ^ ({10{received[131]}} & 10'b0100011100) ^ ({10{received[132]}} & 10'b1000111000) ^ ({10{received[133]}} & 10'b0001111001) ^ ({10{received[134]}} & 10'b0011110010) ^ ({10{received[135]}} & 10'b0111100100) ^ ({10{received[136]}} & 10'b1111001000) ^ ({10{received[137]}} & 10'b1110011001) ^ ({10{received[138]}} & 10'b1100111011) ^ ({10{received[139]}} & 10'b1001111111) ^ ({10{received[140]}} & 10'b0011110111) ^ ({10{received[141]}} & 10'b0111101110) ^ ({10{received[142]}} & 10'b1111011100) ^ ({10{received[143]}} & 10'b1110110001) ^ ({10{received[144]}} & 10'b1101101011) ^ ({10{received[145]}} & 10'b1011011111) ^ ({10{received[146]}} & 10'b0110110111) ^ ({10{received[147]}} & 10'b1101101110) ^ ({10{received[148]}} & 10'b1011010101) ^ ({10{received[149]}} & 10'b0110100011) ^ ({10{received[150]}} & 10'b1101000110) ^ ({10{received[151]}} & 10'b1010000101) ^ ({10{received[152]}} & 10'b0100000011) ^ ({10{received[153]}} & 10'b1000000110) ^ ({10{received[154]}} & 10'b0000000101) ^ ({10{received[155]}} & 10'b0000001010) ^ ({10{received[156]}} & 10'b0000010100) ^ ({10{received[157]}} & 10'b0000101000) ^ ({10{received[158]}} & 10'b0001010000) ^ ({10{received[159]}} & 10'b0010100000) ^ ({10{received[160]}} & 10'b0101000000) ^ ({10{received[161]}} & 10'b1010000000) ^ ({10{received[162]}} & 10'b0100001001) ^ ({10{received[163]}} & 10'b1000010010) ^ ({10{received[164]}} & 10'b0000101101) ^ ({10{received[165]}} & 10'b0001011010) ^ ({10{received[166]}} & 10'b0010110100) ^ ({10{received[167]}} & 10'b0101101000) ^ ({10{received[168]}} & 10'b1011010000) ^ ({10{received[169]}} & 10'b0110101001) ^ ({10{received[170]}} & 10'b1101010010) ^ ({10{received[171]}} & 10'b1010101101) ^ ({10{received[172]}} & 10'b0101010011) ^ ({10{received[173]}} & 10'b1010100110) ^ ({10{received[174]}} & 10'b0101000101) ^ ({10{received[175]}} & 10'b1010001010) ^ ({10{received[176]}} & 10'b0100011101) ^ ({10{received[177]}} & 10'b1000111010) ^ ({10{received[178]}} & 10'b0001111101) ^ ({10{received[179]}} & 10'b0011111010) ^ ({10{received[180]}} & 10'b0111110100) ^ ({10{received[181]}} & 10'b1111101000) ^ ({10{received[182]}} & 10'b1111011001) ^ ({10{received[183]}} & 10'b1110111011) ^ ({10{received[184]}} & 10'b1101111111) ^ ({10{received[185]}} & 10'b1011110111) ^ ({10{received[186]}} & 10'b0111100111) ^ ({10{received[187]}} & 10'b1111001110) ^ ({10{received[188]}} & 10'b1110010101) ^ ({10{received[189]}} & 10'b1100100011) ^ ({10{received[190]}} & 10'b1001001111) ^ ({10{received[191]}} & 10'b0010010111) ^ ({10{received[192]}} & 10'b0100101110) ^ ({10{received[193]}} & 10'b1001011100) ^ ({10{received[194]}} & 10'b0010110001) ^ ({10{received[195]}} & 10'b0101100010) ^ ({10{received[196]}} & 10'b1011000100) ^ ({10{received[197]}} & 10'b0110000001) ^ ({10{received[198]}} & 10'b1100000010) ^ ({10{received[199]}} & 10'b1000001101) ^ ({10{received[200]}} & 10'b0000010011) ^ ({10{received[201]}} & 10'b0000100110) ^ ({10{received[202]}} & 10'b0001001100) ^ ({10{received[203]}} & 10'b0010011000) ^ ({10{received[204]}} & 10'b0100110000) ^ ({10{received[205]}} & 10'b1001100000) ^ ({10{received[206]}} & 10'b0011001001) ^ ({10{received[207]}} & 10'b0110010010) ^ ({10{received[208]}} & 10'b1100100100) ^ ({10{received[209]}} & 10'b1001000001) ^ ({10{received[210]}} & 10'b0010001011) ^ ({10{received[211]}} & 10'b0100010110) ^ ({10{received[212]}} & 10'b1000101100) ^ ({10{received[213]}} & 10'b0001010001) ^ ({10{received[214]}} & 10'b0010100010) ^ ({10{received[215]}} & 10'b0101000100) ^ ({10{received[216]}} & 10'b1010001000) ^ ({10{received[217]}} & 10'b0100011001) ^ ({10{received[218]}} & 10'b1000110010) ^ ({10{received[219]}} & 10'b0001101101) ^ ({10{received[220]}} & 10'b0011011010) ^ ({10{received[221]}} & 10'b0110110100) ^ ({10{received[222]}} & 10'b1101101000) ^ ({10{received[223]}} & 10'b1011011001) ^ ({10{received[224]}} & 10'b0110111011) ^ ({10{received[225]}} & 10'b1101110110) ^ ({10{received[226]}} & 10'b1011100101) ^ ({10{received[227]}} & 10'b0111000011) ^ ({10{received[228]}} & 10'b1110000110) ^ ({10{received[229]}} & 10'b1100000101) ^ ({10{received[230]}} & 10'b1000000011) ^ ({10{received[231]}} & 10'b0000001111) ^ ({10{received[232]}} & 10'b0000011110) ^ ({10{received[233]}} & 10'b0000111100) ^ ({10{received[234]}} & 10'b0001111000) ^ ({10{received[235]}} & 10'b0011110000) ^ ({10{received[236]}} & 10'b0111100000) ^ ({10{received[237]}} & 10'b1111000000) ^ ({10{received[238]}} & 10'b1110001001) ^ ({10{received[239]}} & 10'b1100011011) ^ ({10{received[240]}} & 10'b1000111111) ^ ({10{received[241]}} & 10'b0001110111) ^ ({10{received[242]}} & 10'b0011101110) ^ ({10{received[243]}} & 10'b0111011100) ^ ({10{received[244]}} & 10'b1110111000) ^ ({10{received[245]}} & 10'b1101111001) ^ ({10{received[246]}} & 10'b1011111011) ^ ({10{received[247]}} & 10'b0111111111) ^ ({10{received[248]}} & 10'b1111111110) ^ ({10{received[249]}} & 10'b1111110101) ^ ({10{received[250]}} & 10'b1111100011) ^ ({10{received[251]}} & 10'b1111001111) ^ ({10{received[252]}} & 10'b1110010111) ^ ({10{received[253]}} & 10'b1100100111) ^ ({10{received[254]}} & 10'b1001000111) ^ ({10{received[255]}} & 10'b0010000111) ^ ({10{received[256]}} & 10'b0100001110) ^ ({10{received[257]}} & 10'b1000011100) ^ ({10{received[258]}} & 10'b0000110001) ^ ({10{received[259]}} & 10'b0001100010) ^ ({10{received[260]}} & 10'b0011000100) ^ ({10{received[261]}} & 10'b0110001000) ^ ({10{received[262]}} & 10'b1100010000) ^ ({10{received[263]}} & 10'b1000101001) ^ ({10{received[264]}} & 10'b0001011011) ^ ({10{received[265]}} & 10'b0010110110) ^ ({10{received[266]}} & 10'b0101101100) ^ ({10{received[267]}} & 10'b1011011000) ^ ({10{received[268]}} & 10'b0110111001) ^ ({10{received[269]}} & 10'b1101110010) ^ ({10{received[270]}} & 10'b1011101101) ^ ({10{received[271]}} & 10'b0111010011) ^ ({10{received[272]}} & 10'b1110100110) ^ ({10{received[273]}} & 10'b1101000101) ^ ({10{received[274]}} & 10'b1010000011) ^ ({10{received[275]}} & 10'b0100001111) ^ ({10{received[276]}} & 10'b1000011110) ^ ({10{received[277]}} & 10'b0000110101) ^ ({10{received[278]}} & 10'b0001101010) ^ ({10{received[279]}} & 10'b0011010100) ^ ({10{received[280]}} & 10'b0110101000) ^ ({10{received[281]}} & 10'b1101010000) ^ ({10{received[282]}} & 10'b1010101001) ^ ({10{received[283]}} & 10'b0101011011) ^ ({10{received[284]}} & 10'b1010110110) ^ ({10{received[285]}} & 10'b0101100101) ^ ({10{received[286]}} & 10'b1011001010) ^ ({10{received[287]}} & 10'b0110011101) ^ ({10{received[288]}} & 10'b1100111010) ^ ({10{received[289]}} & 10'b1001111101) ^ ({10{received[290]}} & 10'b0011110011) ^ ({10{received[291]}} & 10'b0111100110) ^ ({10{received[292]}} & 10'b1111001100) ^ ({10{received[293]}} & 10'b1110010001) ^ ({10{received[294]}} & 10'b1100101011) ^ ({10{received[295]}} & 10'b1001011111) ^ ({10{received[296]}} & 10'b0010110111) ^ ({10{received[297]}} & 10'b0101101110) ^ ({10{received[298]}} & 10'b1011011100) ^ ({10{received[299]}} & 10'b0110110001) ^ ({10{received[300]}} & 10'b1101100010) ^ ({10{received[301]}} & 10'b1011001101) ^ ({10{received[302]}} & 10'b0110010011) ^ ({10{received[303]}} & 10'b1100100110) ^ ({10{received[304]}} & 10'b1001000101) ^ ({10{received[305]}} & 10'b0010000011) ^ ({10{received[306]}} & 10'b0100000110) ^ ({10{received[307]}} & 10'b1000001100) ^ ({10{received[308]}} & 10'b0000010001) ^ ({10{received[309]}} & 10'b0000100010) ^ ({10{received[310]}} & 10'b0001000100) ^ ({10{received[311]}} & 10'b0010001000) ^ ({10{received[312]}} & 10'b0100010000) ^ ({10{received[313]}} & 10'b1000100000) ^ ({10{received[314]}} & 10'b0001001001) ^ ({10{received[315]}} & 10'b0010010010) ^ ({10{received[316]}} & 10'b0100100100) ^ ({10{received[317]}} & 10'b1001001000) ^ ({10{received[318]}} & 10'b0010011001) ^ ({10{received[319]}} & 10'b0100110010) ^ ({10{received[320]}} & 10'b1001100100) ^ ({10{received[321]}} & 10'b0011000001) ^ ({10{received[322]}} & 10'b0110000010) ^ ({10{received[323]}} & 10'b1100000100) ^ ({10{received[324]}} & 10'b1000000001) ^ ({10{received[325]}} & 10'b0000001011) ^ ({10{received[326]}} & 10'b0000010110) ^ ({10{received[327]}} & 10'b0000101100) ^ ({10{received[328]}} & 10'b0001011000) ^ ({10{received[329]}} & 10'b0010110000) ^ ({10{received[330]}} & 10'b0101100000) ^ ({10{received[331]}} & 10'b1011000000) ^ ({10{received[332]}} & 10'b0110001001) ^ ({10{received[333]}} & 10'b1100010010) ^ ({10{received[334]}} & 10'b1000101101) ^ ({10{received[335]}} & 10'b0001010011) ^ ({10{received[336]}} & 10'b0010100110) ^ ({10{received[337]}} & 10'b0101001100) ^ ({10{received[338]}} & 10'b1010011000) ^ ({10{received[339]}} & 10'b0100111001) ^ ({10{received[340]}} & 10'b1001110010) ^ ({10{received[341]}} & 10'b0011101101) ^ ({10{received[342]}} & 10'b0111011010) ^ ({10{received[343]}} & 10'b1110110100) ^ ({10{received[344]}} & 10'b1101100001) ^ ({10{received[345]}} & 10'b1011001011) ^ ({10{received[346]}} & 10'b0110011111) ^ ({10{received[347]}} & 10'b1100111110) ^ ({10{received[348]}} & 10'b1001110101) ^ ({10{received[349]}} & 10'b0011100011) ^ ({10{received[350]}} & 10'b0111000110) ^ ({10{received[351]}} & 10'b1110001100) ^ ({10{received[352]}} & 10'b1100010001) ^ ({10{received[353]}} & 10'b1000101011) ^ ({10{received[354]}} & 10'b0001011111) ^ ({10{received[355]}} & 10'b0010111110) ^ ({10{received[356]}} & 10'b0101111100) ^ ({10{received[357]}} & 10'b1011111000) ^ ({10{received[358]}} & 10'b0111111001) ^ ({10{received[359]}} & 10'b1111110010) ^ ({10{received[360]}} & 10'b1111101101) ^ ({10{received[361]}} & 10'b1111010011) ^ ({10{received[362]}} & 10'b1110101111) ^ ({10{received[363]}} & 10'b1101010111) ^ ({10{received[364]}} & 10'b1010100111) ^ ({10{received[365]}} & 10'b0101000111) ^ ({10{received[366]}} & 10'b1010001110) ^ ({10{received[367]}} & 10'b0100010101) ^ ({10{received[368]}} & 10'b1000101010) ^ ({10{received[369]}} & 10'b0001011101) ^ ({10{received[370]}} & 10'b0010111010) ^ ({10{received[371]}} & 10'b0101110100) ^ ({10{received[372]}} & 10'b1011101000) ^ ({10{received[373]}} & 10'b0111011001) ^ ({10{received[374]}} & 10'b1110110010) ^ ({10{received[375]}} & 10'b1101101101) ^ ({10{received[376]}} & 10'b1011010011) ^ ({10{received[377]}} & 10'b0110101111) ^ ({10{received[378]}} & 10'b1101011110) ^ ({10{received[379]}} & 10'b1010110101) ^ ({10{received[380]}} & 10'b0101100011) ^ ({10{received[381]}} & 10'b1011000110) ^ ({10{received[382]}} & 10'b0110000101) ^ ({10{received[383]}} & 10'b1100001010) ^ ({10{received[384]}} & 10'b1000011101) ^ ({10{received[385]}} & 10'b0000110011) ^ ({10{received[386]}} & 10'b0001100110) ^ ({10{received[387]}} & 10'b0011001100) ^ ({10{received[388]}} & 10'b0110011000) ^ ({10{received[389]}} & 10'b1100110000) ^ ({10{received[390]}} & 10'b1001101001) ^ ({10{received[391]}} & 10'b0011011011) ^ ({10{received[392]}} & 10'b0110110110) ^ ({10{received[393]}} & 10'b1101101100) ^ ({10{received[394]}} & 10'b1011010001) ^ ({10{received[395]}} & 10'b0110101011) ^ ({10{received[396]}} & 10'b1101010110) ^ ({10{received[397]}} & 10'b1010100101) ^ ({10{received[398]}} & 10'b0101000011) ^ ({10{received[399]}} & 10'b1010000110) ^ ({10{received[400]}} & 10'b0100000101) ^ ({10{received[401]}} & 10'b1000001010) ^ ({10{received[402]}} & 10'b0000011101) ^ ({10{received[403]}} & 10'b0000111010) ^ ({10{received[404]}} & 10'b0001110100) ^ ({10{received[405]}} & 10'b0011101000) ^ ({10{received[406]}} & 10'b0111010000) ^ ({10{received[407]}} & 10'b1110100000) ^ ({10{received[408]}} & 10'b1101001001) ^ ({10{received[409]}} & 10'b1010011011) ^ ({10{received[410]}} & 10'b0100111111) ^ ({10{received[411]}} & 10'b1001111110) ^ ({10{received[412]}} & 10'b0011110101) ^ ({10{received[413]}} & 10'b0111101010) ^ ({10{received[414]}} & 10'b1111010100) ^ ({10{received[415]}} & 10'b1110100001) ^ ({10{received[416]}} & 10'b1101001011) ^ ({10{received[417]}} & 10'b1010011111) ^ ({10{received[418]}} & 10'b0100110111) ^ ({10{received[419]}} & 10'b1001101110) ^ ({10{received[420]}} & 10'b0011010101) ^ ({10{received[421]}} & 10'b0110101010) ^ ({10{received[422]}} & 10'b1101010100) ^ ({10{received[423]}} & 10'b1010100001) ^ ({10{received[424]}} & 10'b0101001011) ^ ({10{received[425]}} & 10'b1010010110) ^ ({10{received[426]}} & 10'b0100100101) ^ ({10{received[427]}} & 10'b1001001010) ^ ({10{received[428]}} & 10'b0010011101) ^ ({10{received[429]}} & 10'b0100111010) ^ ({10{received[430]}} & 10'b1001110100) ^ ({10{received[431]}} & 10'b0011100001) ^ ({10{received[432]}} & 10'b0111000010) ^ ({10{received[433]}} & 10'b1110000100) ^ ({10{received[434]}} & 10'b1100000001) ^ ({10{received[435]}} & 10'b1000001011) ^ ({10{received[436]}} & 10'b0000011111) ^ ({10{received[437]}} & 10'b0000111110) ^ ({10{received[438]}} & 10'b0001111100) ^ ({10{received[439]}} & 10'b0011111000) ^ ({10{received[440]}} & 10'b0111110000) ^ ({10{received[441]}} & 10'b1111100000) ^ ({10{received[442]}} & 10'b1111001001) ^ ({10{received[443]}} & 10'b1110011011) ^ ({10{received[444]}} & 10'b1100111111) ^ ({10{received[445]}} & 10'b1001110111) ^ ({10{received[446]}} & 10'b0011100111) ^ ({10{received[447]}} & 10'b0111001110) ^ ({10{received[448]}} & 10'b1110011100) ^ ({10{received[449]}} & 10'b1100110001) ^ ({10{received[450]}} & 10'b1001101011) ^ ({10{received[451]}} & 10'b0011011111) ^ ({10{received[452]}} & 10'b0110111110) ^ ({10{received[453]}} & 10'b1101111100) ^ ({10{received[454]}} & 10'b1011110001) ^ ({10{received[455]}} & 10'b0111101011) ^ ({10{received[456]}} & 10'b1111010110) ^ ({10{received[457]}} & 10'b1110100101) ^ ({10{received[458]}} & 10'b1101000011) ^ ({10{received[459]}} & 10'b1010001111) ^ ({10{received[460]}} & 10'b0100010111) ^ ({10{received[461]}} & 10'b1000101110) ^ ({10{received[462]}} & 10'b0001010101) ^ ({10{received[463]}} & 10'b0010101010) ^ ({10{received[464]}} & 10'b0101010100) ^ ({10{received[465]}} & 10'b1010101000) ^ ({10{received[466]}} & 10'b0101011001) ^ ({10{received[467]}} & 10'b1010110010) ^ ({10{received[468]}} & 10'b0101101101) ^ ({10{received[469]}} & 10'b1011011010) ^ ({10{received[470]}} & 10'b0110111101) ^ ({10{received[471]}} & 10'b1101111010) ^ ({10{received[472]}} & 10'b1011111101) ^ ({10{received[473]}} & 10'b0111110011) ^ ({10{received[474]}} & 10'b1111100110) ^ ({10{received[475]}} & 10'b1111000101) ^ ({10{received[476]}} & 10'b1110000011) ^ ({10{received[477]}} & 10'b1100001111) ^ ({10{received[478]}} & 10'b1000010111) ^ ({10{received[479]}} & 10'b0000100111) ^ ({10{received[480]}} & 10'b0001001110) ^ ({10{received[481]}} & 10'b0010011100) ^ ({10{received[482]}} & 10'b0100111000) ^ ({10{received[483]}} & 10'b1001110000) ^ ({10{received[484]}} & 10'b0011101001) ^ ({10{received[485]}} & 10'b0111010010) ^ ({10{received[486]}} & 10'b1110100100) ^ ({10{received[487]}} & 10'b1101000001) ^ ({10{received[488]}} & 10'b1010001011) ^ ({10{received[489]}} & 10'b0100011111) ^ ({10{received[490]}} & 10'b1000111110) ^ ({10{received[491]}} & 10'b0001110101) ^ ({10{received[492]}} & 10'b0011101010) ^ ({10{received[493]}} & 10'b0111010100) ^ ({10{received[494]}} & 10'b1110101000) ^ ({10{received[495]}} & 10'b1101011001) ^ ({10{received[496]}} & 10'b1010111011) ^ ({10{received[497]}} & 10'b0101111111) ^ ({10{received[498]}} & 10'b1011111110) ^ ({10{received[499]}} & 10'b0111110101) ^ ({10{received[500]}} & 10'b1111101010) ^ ({10{received[501]}} & 10'b1111011101) ^ ({10{received[502]}} & 10'b1110110011) ^ ({10{received[503]}} & 10'b1101101111) ^ ({10{received[504]}} & 10'b1011010111) ^ ({10{received[505]}} & 10'b0110100111) ^ ({10{received[506]}} & 10'b1101001110) ^ ({10{received[507]}} & 10'b1010010101) ^ ({10{received[508]}} & 10'b0100100011) ^ ({10{received[509]}} & 10'b1001000110) ^ ({10{received[510]}} & 10'b0010000101) ^ ({10{received[511]}} & 10'b0100001010) ^ ({10{received[512]}} & 10'b1000010100) ^ ({10{received[513]}} & 10'b0000100001) ^ ({10{received[514]}} & 10'b0001000010) ^ ({10{received[515]}} & 10'b0010000100) ^ ({10{received[516]}} & 10'b0100001000) ^ ({10{received[517]}} & 10'b1000010000) ^ ({10{received[518]}} & 10'b0000101001) ^ ({10{received[519]}} & 10'b0001010010) ^ ({10{received[520]}} & 10'b0010100100) ^ ({10{received[521]}} & 10'b0101001000) ^ ({10{received[522]}} & 10'b1010010000) ^ ({10{received[523]}} & 10'b0100101001) ^ ({10{received[524]}} & 10'b1001010010) ^ ({10{received[525]}} & 10'b0010101101) ^ ({10{received[526]}} & 10'b0101011010) ^ ({10{received[527]}} & 10'b1010110100) ^ ({10{received[528]}} & 10'b0101100001) ^ ({10{received[529]}} & 10'b1011000010) ^ ({10{received[530]}} & 10'b0110001101) ^ ({10{received[531]}} & 10'b1100011010) ^ ({10{received[532]}} & 10'b1000111101) ^ ({10{received[533]}} & 10'b0001110011) ^ ({10{received[534]}} & 10'b0011100110) ^ ({10{received[535]}} & 10'b0111001100) ^ ({10{received[536]}} & 10'b1110011000) ^ ({10{received[537]}} & 10'b1100111001) ^ ({10{received[538]}} & 10'b1001111011) ^ ({10{received[539]}} & 10'b0011111111) ^ ({10{received[540]}} & 10'b0111111110) ^ ({10{received[541]}} & 10'b1111111100);
  assign syndrome2 = ({10{received[0]}} & 10'b0000000001) ^ 
  ({10{received[1]}} & 10'b0000000100) ^ ({10{received[2]}} & 10'b0000010000) ^ ({10{received[3]}} & 10'b0001000000) ^ ({10{received[4]}} & 10'b0100000000) ^ ({10{received[5]}} & 10'b0000001001) ^ ({10{received[6]}} & 10'b0000100100) ^ ({10{received[7]}} & 10'b0010010000) ^ ({10{received[8]}} & 10'b1001000000) ^ ({10{received[9]}} & 10'b0100010010) ^ ({10{received[10]}} & 10'b0001000001) ^ ({10{received[11]}} & 10'b0100000100) ^ ({10{received[12]}} & 10'b0000011001) ^ ({10{received[13]}} & 10'b0001100100) ^ ({10{received[14]}} & 10'b0110010000) ^ ({10{received[15]}} & 10'b1001001001) ^ ({10{received[16]}} & 10'b0100110110) ^ ({10{received[17]}} & 10'b0011010001) ^ ({10{received[18]}} & 10'b1101000100) ^ ({10{received[19]}} & 10'b0100001011) ^ ({10{received[20]}} & 10'b0000100101) ^ ({10{received[21]}} & 10'b0010010100) ^ ({10{received[22]}} & 10'b1001010000) ^ ({10{received[23]}} & 10'b0101010010) ^ ({10{received[24]}} & 10'b0101000001) ^ ({10{received[25]}} & 10'b0100001101) ^ ({10{received[26]}} & 10'b0000111101) ^ ({10{received[27]}} & 10'b0011110100) ^ ({10{received[28]}} & 10'b1111010000) ^ ({10{received[29]}} & 10'b1101011011) ^ ({10{received[30]}} & 10'b0101110111) ^ ({10{received[31]}} & 10'b0111010101) ^ ({10{received[32]}} & 10'b1101011101) ^ ({10{received[33]}} & 10'b0101101111) ^ ({10{received[34]}} & 10'b0110110101) ^ ({10{received[35]}} & 10'b1011011101) ^ ({10{received[36]}} & 10'b1101100110) ^ ({10{received[37]}} & 10'b0110000011) ^ ({10{received[38]}} & 10'b1000000101) ^ ({10{received[39]}} & 10'b0000000110) ^ ({10{received[40]}} & 10'b0000011000) ^ ({10{received[41]}} & 10'b0001100000) ^ ({10{received[42]}} & 10'b0110000000) ^ ({10{received[43]}} & 10'b1000001001) ^ ({10{received[44]}} & 10'b0000110110) ^ ({10{received[45]}} & 10'b0011011000) ^ ({10{received[46]}} & 10'b1101100000) ^ ({10{received[47]}} & 10'b0110011011) ^ ({10{received[48]}} & 10'b1001100101) ^ ({10{received[49]}} & 10'b0110000110) ^ ({10{received[50]}} & 10'b1000010001) ^ ({10{received[51]}} & 10'b0001010110) ^ ({10{received[52]}} & 10'b0101011000) ^ ({10{received[53]}} & 10'b0101101001) ^ ({10{received[54]}} & 10'b0110101101) ^ ({10{received[55]}} & 10'b1010111101) ^ ({10{received[56]}} & 10'b1011100110) ^ ({10{received[57]}} & 10'b1110001010) ^ ({10{received[58]}} & 10'b1000110011) ^ ({10{received[59]}} & 10'b0011011110) ^ ({10{received[60]}} & 10'b1101111000) ^ ({10{received[61]}} & 10'b0111111011) ^ ({10{received[62]}} & 10'b1111100101) ^ ({10{received[63]}} & 10'b1110001111) ^ ({10{received[64]}} & 10'b1000100111) ^ ({10{received[65]}} & 10'b0010001110) ^ ({10{received[66]}} & 10'b1000111000) ^ ({10{received[67]}} & 10'b0011110010) ^ ({10{received[68]}} & 10'b1111001000) ^ ({10{received[69]}} & 10'b1100111011) ^ ({10{received[70]}} & 10'b0011110111) ^ ({10{received[71]}} & 10'b1111011100) ^ ({10{received[72]}} & 10'b1101101011) ^ ({10{received[73]}} & 10'b0110110111) ^ ({10{received[74]}} & 10'b1011010101) ^ ({10{received[75]}} & 10'b1101000110) ^ ({10{received[76]}} & 10'b0100000011) ^ ({10{received[77]}} & 10'b0000000101) ^ ({10{received[78]}} & 10'b0000010100) ^ ({10{received[79]}} & 10'b0001010000) ^ ({10{received[80]}} & 10'b0101000000) ^ ({10{received[81]}} & 10'b0100001001) ^ ({10{received[82]}} & 10'b0000101101) ^ ({10{received[83]}} & 10'b0010110100) ^ ({10{received[84]}} & 10'b1011010000) ^ ({10{received[85]}} & 10'b1101010010) ^ ({10{received[86]}} & 10'b0101010011) ^ ({10{received[87]}} & 10'b0101000101) ^ ({10{received[88]}} & 10'b0100011101) ^ ({10{received[89]}} & 10'b0001111101) ^ ({10{received[90]}} & 10'b0111110100) ^ ({10{received[91]}} & 10'b1111011001) ^ ({10{received[92]}} & 10'b1101111111) ^ ({10{received[93]}} & 10'b0111100111) ^ ({10{received[94]}} & 10'b1110010101) ^ ({10{received[95]}} & 10'b1001001111) ^ ({10{received[96]}} & 10'b0100101110) ^ ({10{received[97]}} & 10'b0010110001) ^ ({10{received[98]}} & 10'b1011000100) ^ ({10{received[99]}} & 10'b1100000010) ^ ({10{received[100]}} & 10'b0000010011) ^ ({10{received[101]}} & 10'b0001001100) ^ ({10{received[102]}} & 10'b0100110000) ^ ({10{received[103]}} & 10'b0011001001) ^ ({10{received[104]}} & 10'b1100100100) ^ ({10{received[105]}} & 10'b0010001011) ^ ({10{received[106]}} & 10'b1000101100) ^ ({10{received[107]}} & 10'b0010100010) ^ ({10{received[108]}} & 10'b1010001000) ^ ({10{received[109]}} & 10'b1000110010) ^ ({10{received[110]}} & 10'b0011011010) ^ ({10{received[111]}} & 10'b1101101000) ^ ({10{received[112]}} & 10'b0110111011) ^ ({10{received[113]}} & 10'b1011100101) ^ ({10{received[114]}} & 10'b1110000110) ^ ({10{received[115]}} & 10'b1000000011) ^ ({10{received[116]}} & 10'b0000011110) ^ ({10{received[117]}} & 10'b0001111000) ^ ({10{received[118]}} & 10'b0111100000) ^ ({10{received[119]}} & 10'b1110001001) ^ ({10{received[120]}} & 10'b1000111111) ^ ({10{received[121]}} & 10'b0011101110) ^ ({10{received[122]}} & 10'b1110111000) ^ ({10{received[123]}} & 10'b1011111011) ^ ({10{received[124]}} & 10'b1111111110) ^ ({10{received[125]}} & 10'b1111100011) ^ ({10{received[126]}} & 10'b1110010111) ^ ({10{received[127]}} & 10'b1001000111) ^ ({10{received[128]}} & 10'b0100001110) ^ ({10{received[129]}} & 10'b0000110001) ^ ({10{received[130]}} & 10'b0011000100) ^ ({10{received[131]}} & 10'b1100010000) ^ ({10{received[132]}} & 10'b0001011011) ^ ({10{received[133]}} & 10'b0101101100) ^ ({10{received[134]}} & 10'b0110111001) ^ ({10{received[135]}} & 10'b1011101101) ^ ({10{received[136]}} & 10'b1110100110) ^ ({10{received[137]}} & 10'b1010000011) ^ ({10{received[138]}} & 10'b1000011110) ^ ({10{received[139]}} & 10'b0001101010) ^ ({10{received[140]}} & 10'b0110101000) ^ ({10{received[141]}} & 10'b1010101001) ^ ({10{received[142]}} & 10'b1010110110) ^ ({10{received[143]}} & 10'b1011001010) ^ ({10{received[144]}} & 10'b1100111010) ^ ({10{received[145]}} & 10'b0011110011) ^ ({10{received[146]}} & 10'b1111001100) ^ ({10{received[147]}} & 10'b1100101011) ^ ({10{received[148]}} & 10'b0010110111) ^ ({10{received[149]}} & 10'b1011011100) ^ ({10{received[150]}} & 10'b1101100010) ^ ({10{received[151]}} & 10'b0110010011) ^ ({10{received[152]}} & 10'b1001000101) ^ ({10{received[153]}} & 10'b0100000110) ^ ({10{received[154]}} & 10'b0000010001) ^ ({10{received[155]}} & 10'b0001000100) ^ ({10{received[156]}} & 10'b0100010000) ^ ({10{received[157]}} & 10'b0001001001) ^ ({10{received[158]}} & 10'b0100100100) ^ ({10{received[159]}} & 10'b0010011001) ^ ({10{received[160]}} & 10'b1001100100) ^ ({10{received[161]}} & 10'b0110000010) ^ ({10{received[162]}} & 10'b1000000001) ^ ({10{received[163]}} & 10'b0000010110) ^ ({10{received[164]}} & 10'b0001011000) ^ ({10{received[165]}} & 10'b0101100000) ^ ({10{received[166]}} & 10'b0110001001) ^ ({10{received[167]}} & 10'b1000101101) ^ ({10{received[168]}} & 10'b0010100110) ^ ({10{received[169]}} & 10'b1010011000) ^ ({10{received[170]}} & 10'b1001110010) ^ ({10{received[171]}} & 10'b0111011010) ^ ({10{received[172]}} & 10'b1101100001) ^ ({10{received[173]}} & 10'b0110011111) ^ ({10{received[174]}} & 10'b1001110101) ^ ({10{received[175]}} & 10'b0111000110) ^ ({10{received[176]}} & 10'b1100010001) ^ ({10{received[177]}} & 10'b0001011111) ^ ({10{received[178]}} & 10'b0101111100) ^ ({10{received[179]}} & 10'b0111111001) ^ ({10{received[180]}} & 10'b1111101101) ^ ({10{received[181]}} & 10'b1110101111) ^ ({10{received[182]}} & 10'b1010100111) ^ ({10{received[183]}} & 10'b1010001110) ^ ({10{received[184]}} & 10'b1000101010) ^ ({10{received[185]}} & 10'b0010111010) ^ ({10{received[186]}} & 10'b1011101000) ^ ({10{received[187]}} & 10'b1110110010) ^ ({10{received[188]}} & 10'b1011010011) ^ ({10{received[189]}} & 10'b1101011110) ^ ({10{received[190]}} & 10'b0101100011) ^ ({10{received[191]}} & 10'b0110000101) ^ ({10{received[192]}} & 10'b1000011101) ^ ({10{received[193]}} & 10'b0001100110) ^ ({10{received[194]}} & 10'b0110011000) ^ ({10{received[195]}} & 10'b1001101001) ^ ({10{received[196]}} & 10'b0110110110) ^ ({10{received[197]}} & 10'b1011010001) ^ ({10{received[198]}} & 10'b1101010110) ^ ({10{received[199]}} & 10'b0101000011) ^ ({10{received[200]}} & 10'b0100000101) ^ ({10{received[201]}} & 10'b0000011101) ^ ({10{received[202]}} & 10'b0001110100) ^ ({10{received[203]}} & 10'b0111010000) ^ ({10{received[204]}} & 10'b1101001001) ^ ({10{received[205]}} & 10'b0100111111) ^ ({10{received[206]}} & 10'b0011110101) ^ ({10{received[207]}} & 10'b1111010100) ^ ({10{received[208]}} & 10'b1101001011) ^ ({10{received[209]}} & 10'b0100110111) ^ ({10{received[210]}} & 10'b0011010101) ^ ({10{received[211]}} & 10'b1101010100) ^ ({10{received[212]}} & 10'b0101001011) ^ ({10{received[213]}} & 10'b0100100101) ^ ({10{received[214]}} & 10'b0010011101) ^ ({10{received[215]}} & 10'b1001110100) ^ ({10{received[216]}} & 10'b0111000010) ^ ({10{received[217]}} & 10'b1100000001) ^ ({10{received[218]}} & 10'b0000011111) ^ ({10{received[219]}} & 10'b0001111100) ^ ({10{received[220]}} & 10'b0111110000) ^ ({10{received[221]}} & 10'b1111001001) ^ ({10{received[222]}} & 10'b1100111111) ^ ({10{received[223]}} & 10'b0011100111) ^ ({10{received[224]}} & 10'b1110011100) ^ ({10{received[225]}} & 10'b1001101011) ^ ({10{received[226]}} & 10'b0110111110) ^ ({10{received[227]}} & 10'b1011110001) ^ ({10{received[228]}} & 10'b1111010110) ^ ({10{received[229]}} & 10'b1101000011) ^ ({10{received[230]}} & 10'b0100010111) ^ ({10{received[231]}} & 10'b0001010101) ^ ({10{received[232]}} & 10'b0101010100) ^ ({10{received[233]}} & 10'b0101011001) ^ ({10{received[234]}} & 10'b0101101101) ^ ({10{received[235]}} & 10'b0110111101) ^ ({10{received[236]}} & 10'b1011111101) ^ ({10{received[237]}} & 10'b1111100110) ^ ({10{received[238]}} & 10'b1110000011) ^ ({10{received[239]}} & 10'b1000010111) ^ ({10{received[240]}} & 10'b0001001110) ^ ({10{received[241]}} & 10'b0100111000) ^ ({10{received[242]}} & 10'b0011101001) ^ ({10{received[243]}} & 10'b1110100100) ^ ({10{received[244]}} & 10'b1010001011) ^ ({10{received[245]}} & 10'b1000111110) ^ ({10{received[246]}} & 10'b0011101010) ^ ({10{received[247]}} & 10'b1110101000) ^ ({10{received[248]}} & 10'b1010111011) ^ ({10{received[249]}} & 10'b1011111110) ^ ({10{received[250]}} & 10'b1111101010) ^ ({10{received[251]}} & 10'b1110110011) ^ ({10{received[252]}} & 10'b1011010111) ^ ({10{received[253]}} & 10'b1101001110) ^ ({10{received[254]}} & 10'b0100100011) ^ ({10{received[255]}} & 10'b0010000101) ^ ({10{received[256]}} & 10'b1000010100) ^ ({10{received[257]}} & 10'b0001000010) ^ ({10{received[258]}} & 10'b0100001000) ^ ({10{received[259]}} & 10'b0000101001) ^ ({10{received[260]}} & 10'b0010100100) ^ ({10{received[261]}} & 10'b1010010000) ^ ({10{received[262]}} & 10'b1001010010) ^ ({10{received[263]}} & 10'b0101011010) ^ ({10{received[264]}} & 10'b0101100001) ^ ({10{received[265]}} & 10'b0110001101) ^ ({10{received[266]}} & 10'b1000111101) ^ ({10{received[267]}} & 10'b0011100110) ^ ({10{received[268]}} & 10'b1110011000) ^ ({10{received[269]}} & 10'b1001111011) ^ ({10{received[270]}} & 10'b0111111110) ^ ({10{received[271]}} & 10'b1111110001) ^ ({10{received[272]}} & 10'b1111011111) ^ ({10{received[273]}} & 10'b1101100111) ^ ({10{received[274]}} & 10'b0110000111) ^ ({10{received[275]}} & 10'b1000010101) ^ ({10{received[276]}} & 10'b0001000110) ^ ({10{received[277]}} & 10'b0100011000) ^ ({10{received[278]}} & 10'b0001101001) ^ ({10{received[279]}} & 10'b0110100100) ^ ({10{received[280]}} & 10'b1010011001) ^ ({10{received[281]}} & 10'b1001110110) ^ ({10{received[282]}} & 10'b0111001010) ^ ({10{received[283]}} & 10'b1100100001) ^ ({10{received[284]}} & 10'b0010011111) ^ ({10{received[285]}} & 10'b1001111100) ^ ({10{received[286]}} & 10'b0111100010) ^ ({10{received[287]}} & 10'b1110000001) ^ ({10{received[288]}} & 10'b1000011111) ^ ({10{received[289]}} & 10'b0001101110) ^ ({10{received[290]}} & 10'b0110111000) ^ ({10{received[291]}} & 10'b1011101001) ^ ({10{received[292]}} & 10'b1110110110) ^ ({10{received[293]}} & 10'b1011000011) ^ ({10{received[294]}} & 10'b1100011110) ^ ({10{received[295]}} & 10'b0001100011) ^ ({10{received[296]}} & 10'b0110001100) ^ ({10{received[297]}} & 10'b1000111001) ^ ({10{received[298]}} & 10'b0011110110) ^ ({10{received[299]}} & 10'b1111011000) ^ ({10{received[300]}} & 10'b1101111011) ^ ({10{received[301]}} & 10'b0111110111) ^ ({10{received[302]}} & 10'b1111010101) ^ ({10{received[303]}} & 10'b1101001111) ^ ({10{received[304]}} & 10'b0100100111) ^ ({10{received[305]}} & 10'b0010010101) ^ ({10{received[306]}} & 10'b1001010100) ^ ({10{received[307]}} & 10'b0101000010) ^ ({10{received[308]}} & 10'b0100000001) ^ ({10{received[309]}} & 10'b0000001101) ^ ({10{received[310]}} & 10'b0000110100) ^ ({10{received[311]}} & 10'b0011010000) ^ ({10{received[312]}} & 10'b1101000000) ^ ({10{received[313]}} & 10'b0100011011) ^ ({10{received[314]}} & 10'b0001100101) ^ ({10{received[315]}} & 10'b0110010100) ^ ({10{received[316]}} & 10'b1001011001) ^ ({10{received[317]}} & 10'b0101110110) ^ ({10{received[318]}} & 10'b0111010001) ^ ({10{received[319]}} & 10'b1101001101) ^ ({10{received[320]}} & 10'b0100101111) ^ ({10{received[321]}} & 10'b0010110101) ^ ({10{received[322]}} & 10'b1011010100) ^ ({10{received[323]}} & 10'b1101000010) ^ ({10{received[324]}} & 10'b0100010011) ^ ({10{received[325]}} & 10'b0001000101) ^ ({10{received[326]}} & 10'b0100010100) ^ ({10{received[327]}} & 10'b0001011001) ^ ({10{received[328]}} & 10'b0101100100) ^ ({10{received[329]}} & 10'b0110011001) ^ ({10{received[330]}} & 10'b1001101101) ^ ({10{received[331]}} & 10'b0110100110) ^ ({10{received[332]}} & 10'b1010010001) ^ ({10{received[333]}} & 10'b1001010110) ^ ({10{received[334]}} & 10'b0101001010) ^ ({10{received[335]}} & 10'b0100100001) ^ ({10{received[336]}} & 10'b0010001101) ^ ({10{received[337]}} & 10'b1000110100) ^ ({10{received[338]}} & 10'b0011000010) ^ ({10{received[339]}} & 10'b1100001000) ^ ({10{received[340]}} & 10'b0000111011) ^ ({10{received[341]}} & 10'b0011101100) ^ ({10{received[342]}} & 10'b1110110000) ^ ({10{received[343]}} & 10'b1011011011) ^ ({10{received[344]}} & 10'b1101111110) ^ ({10{received[345]}} & 10'b0111100011) ^ ({10{received[346]}} & 10'b1110000101) ^ ({10{received[347]}} & 10'b1000001111) ^ ({10{received[348]}} & 10'b0000101110) ^ ({10{received[349]}} & 10'b0010111000) ^ ({10{received[350]}} & 10'b1011100000) ^ ({10{received[351]}} & 10'b1110010010) ^ ({10{received[352]}} & 10'b1001010011) ^ ({10{received[353]}} & 10'b0101011110) ^ ({10{received[354]}} & 10'b0101110001) ^ ({10{received[355]}} & 10'b0111001101) ^ ({10{received[356]}} & 10'b1100111101) ^ ({10{received[357]}} & 10'b0011101111) ^ ({10{received[358]}} & 10'b1110111100) ^ ({10{received[359]}} & 10'b1011101011) ^ ({10{received[360]}} & 10'b1110111110) ^ ({10{received[361]}} & 10'b1011100011) ^ ({10{received[362]}} & 10'b1110011110) ^ ({10{received[363]}} & 10'b1001100011) ^ ({10{received[364]}} & 10'b0110011110) ^ ({10{received[365]}} & 10'b1001110001) ^ ({10{received[366]}} & 10'b0111010110) ^ ({10{received[367]}} & 10'b1101010001) ^ ({10{received[368]}} & 10'b0101011111) ^ ({10{received[369]}} & 10'b0101110101) ^ ({10{received[370]}} & 10'b0111011101) ^ ({10{received[371]}} & 10'b1101111101) ^ ({10{received[372]}} & 10'b0111101111) ^ ({10{received[373]}} & 10'b1110110101) ^ ({10{received[374]}} & 10'b1011001111) ^ ({10{received[375]}} & 10'b1100101110) ^ ({10{received[376]}} & 10'b0010100011) ^ ({10{received[377]}} & 10'b1010001100) ^ ({10{received[378]}} & 10'b1000100010) ^ ({10{received[379]}} & 10'b0010011010) ^ ({10{received[380]}} & 10'b1001101000) ^ ({10{received[381]}} & 10'b0110110010) ^ ({10{received[382]}} & 10'b1011000001) ^ ({10{received[383]}} & 10'b1100010110) ^ ({10{received[384]}} & 10'b0001000011) ^ ({10{received[385]}} & 10'b0100001100) ^ ({10{received[386]}} & 10'b0000111001) ^ ({10{received[387]}} & 10'b0011100100) ^ ({10{received[388]}} & 10'b1110010000) ^ ({10{received[389]}} & 10'b1001011011) ^ ({10{received[390]}} & 10'b0101111110) ^ ({10{received[391]}} & 10'b0111110001) ^ ({10{received[392]}} & 10'b1111001101) ^ ({10{received[393]}} & 10'b1100101111) ^ ({10{received[394]}} & 10'b0010100111) ^ ({10{received[395]}} & 10'b1010011100) ^ ({10{received[396]}} & 10'b1001100010) ^ ({10{received[397]}} & 10'b0110011010) ^ ({10{received[398]}} & 10'b1001100001) ^ ({10{received[399]}} & 10'b0110010110) ^ ({10{received[400]}} & 10'b1001010001) ^ ({10{received[401]}} & 10'b0101010110) ^ ({10{received[402]}} & 10'b0101010001) ^ ({10{received[403]}} & 10'b0101001101) ^ ({10{received[404]}} & 10'b0100111101) ^ ({10{received[405]}} & 10'b0011111101) ^ ({10{received[406]}} & 10'b1111110100) ^ ({10{received[407]}} & 10'b1111001011) ^ ({10{received[408]}} & 10'b1100110111) ^ ({10{received[409]}} & 10'b0011000111) ^ ({10{received[410]}} & 10'b1100011100) ^ ({10{received[411]}} & 10'b0001101011) ^ ({10{received[412]}} & 10'b0110101100) ^ ({10{received[413]}} & 10'b1010111001) ^ ({10{received[414]}} & 10'b1011110110) ^ ({10{received[415]}} & 10'b1111001010) ^ ({10{received[416]}} & 10'b1100110011) ^ ({10{received[417]}} & 10'b0011010111) ^ ({10{received[418]}} & 10'b1101011100) ^ ({10{received[419]}} & 10'b0101101011) ^ ({10{received[420]}} & 10'b0110100101) ^ ({10{received[421]}} & 10'b1010011101) ^ ({10{received[422]}} & 10'b1001100110) ^ ({10{received[423]}} & 10'b0110001010) ^ ({10{received[424]}} & 10'b1000100001) ^ ({10{received[425]}} & 10'b0010010110) ^ ({10{received[426]}} & 10'b1001011000) ^ ({10{received[427]}} & 10'b0101110010) ^ ({10{received[428]}} & 10'b0111000001) ^ ({10{received[429]}} & 10'b1100001101) ^ ({10{received[430]}} & 10'b0000101111) ^ ({10{received[431]}} & 10'b0010111100) ^ ({10{received[432]}} & 10'b1011110000) ^ ({10{received[433]}} & 10'b1111010010) ^ ({10{received[434]}} & 10'b1101010011) ^ ({10{received[435]}} & 10'b0101010111) ^ ({10{received[436]}} & 10'b0101010101) ^ ({10{received[437]}} & 10'b0101011101) ^ ({10{received[438]}} & 10'b0101111101) ^ ({10{received[439]}} & 10'b0111111101) ^ ({10{received[440]}} & 10'b1111111101) ^ ({10{received[441]}} & 10'b1111101111) ^ ({10{received[442]}} & 10'b1110100111) ^ ({10{received[443]}} & 10'b1010000111) ^ ({10{received[444]}} & 10'b1000001110) ^ ({10{received[445]}} & 10'b0000101010) ^ ({10{received[446]}} & 10'b0010101000) ^ ({10{received[447]}} & 10'b1010100000) ^ ({10{received[448]}} & 10'b1010010010) ^ ({10{received[449]}} & 10'b1001011010) ^ ({10{received[450]}} & 10'b0101111010) ^ ({10{received[451]}} & 10'b0111100001) ^ ({10{received[452]}} & 10'b1110001101) ^ ({10{received[453]}} & 10'b1000101111) ^ ({10{received[454]}} & 10'b0010101110) ^ ({10{received[455]}} & 10'b1010111000) ^ ({10{received[456]}} & 10'b1011110010) ^ ({10{received[457]}} & 10'b1111011010) ^ ({10{received[458]}} & 10'b1101110011) ^ ({10{received[459]}} & 10'b0111010111) ^ ({10{received[460]}} & 10'b1101010101) ^ ({10{received[461]}} & 10'b0101001111) ^ ({10{received[462]}} & 10'b0100110101) ^ ({10{received[463]}} & 10'b0011011101) ^ ({10{received[464]}} & 10'b1101110100) ^ ({10{received[465]}} & 10'b0111001011) ^ ({10{received[466]}} & 10'b1100100101) ^ ({10{received[467]}} & 10'b0010001111) ^ ({10{received[468]}} & 10'b1000111100) ^ ({10{received[469]}} & 10'b0011100010) ^ ({10{received[470]}} & 10'b1110001000) ^ ({10{received[471]}} & 10'b1000111011) ^ ({10{received[472]}} & 10'b0011111110) ^ ({10{received[473]}} & 10'b1111111000) ^ ({10{received[474]}} & 10'b1111111011) ^ ({10{received[475]}} & 10'b1111110111) ^ ({10{received[476]}} & 10'b1111000111) ^ ({10{received[477]}} & 10'b1100000111) ^ ({10{received[478]}} & 10'b0000000111) ^ ({10{received[479]}} & 10'b0000011100) ^ ({10{received[480]}} & 10'b0001110000) ^ ({10{received[481]}} & 10'b0111000000) ^ ({10{received[482]}} & 10'b1100001001) ^ ({10{received[483]}} & 10'b0000111111) ^ ({10{received[484]}} & 10'b0011111100) ^ ({10{received[485]}} & 10'b1111110000) ^ ({10{received[486]}} & 10'b1111011011) ^ ({10{received[487]}} & 10'b1101110111) ^ ({10{received[488]}} & 10'b0111000111) ^ ({10{received[489]}} & 10'b1100010101) ^ ({10{received[490]}} & 10'b0001001111) ^ ({10{received[491]}} & 10'b0100111100) ^ ({10{received[492]}} & 10'b0011111001) ^ ({10{received[493]}} & 10'b1111100100) ^ ({10{received[494]}} & 10'b1110001011) ^ ({10{received[495]}} & 10'b1000110111) ^ ({10{received[496]}} & 10'b0011001110) ^ ({10{received[497]}} & 10'b1100111000) ^ ({10{received[498]}} & 10'b0011111011) ^ ({10{received[499]}} & 10'b1111101100) ^ ({10{received[500]}} & 10'b1110101011) ^ ({10{received[501]}} & 10'b1010110111) ^ ({10{received[502]}} & 10'b1011001110) ^ ({10{received[503]}} & 10'b1100101010) ^ ({10{received[504]}} & 10'b0010110011) ^ ({10{received[505]}} & 10'b1011001100) ^ ({10{received[506]}} & 10'b1100100010) ^ ({10{received[507]}} & 10'b0010010011) ^ ({10{received[508]}} & 10'b1001001100) ^ ({10{received[509]}} & 10'b0100100010) ^ ({10{received[510]}} & 10'b0010000001) ^ ({10{received[511]}} & 10'b1000000100) ^ ({10{received[512]}} & 10'b0000000010) ^ ({10{received[513]}} & 10'b0000001000) ^ ({10{received[514]}} & 10'b0000100000) ^ ({10{received[515]}} & 10'b0010000000) ^ ({10{received[516]}} & 10'b1000000000) ^ ({10{received[517]}} & 10'b0000010010) ^ ({10{received[518]}} & 10'b0001001000) ^ ({10{received[519]}} & 10'b0100100000) ^ ({10{received[520]}} & 10'b0010001001) ^ ({10{received[521]}} & 10'b1000100100) ^ ({10{received[522]}} & 10'b0010000010) ^ ({10{received[523]}} & 10'b1000001000) ^ ({10{received[524]}} & 10'b0000110010) ^ ({10{received[525]}} & 10'b0011001000) ^ ({10{received[526]}} & 10'b1100100000) ^ ({10{received[527]}} & 10'b0010011011) ^ ({10{received[528]}} & 10'b1001101100) ^ ({10{received[529]}} & 10'b0110100010) ^ ({10{received[530]}} & 10'b1010000001) ^ ({10{received[531]}} & 10'b1000010110) ^ ({10{received[532]}} & 10'b0001001010) ^ ({10{received[533]}} & 10'b0100101000) ^ ({10{received[534]}} & 10'b0010101001) ^ ({10{received[535]}} & 10'b1010100100) ^ ({10{received[536]}} & 10'b1010000010) ^ ({10{received[537]}} & 10'b1000011010) ^ ({10{received[538]}} & 10'b0001111010) ^ ({10{received[539]}} & 10'b0111101000) ^ ({10{received[540]}} & 10'b1110101001) ^ ({10{received[541]}} & 10'b1010111111);
  assign syndrome3 = ({10{received[0]}} & 10'b0000000001) ^ 
  ({10{received[1]}} & 10'b0000001000) ^ ({10{received[2]}} & 10'b0001000000) ^ ({10{received[3]}} & 10'b1000000000) ^ ({10{received[4]}} & 10'b0000100100) ^ ({10{received[5]}} & 10'b0100100000) ^ ({10{received[6]}} & 10'b0100010010) ^ ({10{received[7]}} & 10'b0010000010) ^ ({10{received[8]}} & 10'b0000011001) ^ ({10{received[9]}} & 10'b0011001000) ^ ({10{received[10]}} & 10'b1001001001) ^ ({10{received[11]}} & 10'b1001101100) ^ ({10{received[12]}} & 10'b1101000100) ^ ({10{received[13]}} & 10'b1000010110) ^ ({10{received[14]}} & 10'b0010010100) ^ ({10{received[15]}} & 10'b0010101001) ^ ({10{received[16]}} & 10'b0101000001) ^ ({10{received[17]}} & 10'b1000011010) ^ ({10{received[18]}} & 10'b0011110100) ^ ({10{received[19]}} & 10'b1110101001) ^ ({10{received[20]}} & 10'b0101110111) ^ ({10{received[21]}} & 10'b1110101010) ^ ({10{received[22]}} & 10'b0101101111) ^ ({10{received[23]}} & 10'b1101101010) ^ ({10{received[24]}} & 10'b1101100110) ^ ({10{received[25]}} & 10'b1100000110) ^ ({10{received[26]}} & 10'b0000000110) ^ ({10{received[27]}} & 10'b0000110000) ^ ({10{received[28]}} & 10'b0110000000) ^ ({10{received[29]}} & 10'b0000011011) ^ ({10{received[30]}} & 10'b0011011000) ^ ({10{received[31]}} & 10'b1011001001) ^ ({10{received[32]}} & 10'b1001100101) ^ ({10{received[33]}} & 10'b1100001100) ^ ({10{received[34]}} & 10'b0001010110) ^ ({10{received[35]}} & 10'b1010110000) ^ ({10{received[36]}} & 10'b0110101101) ^ ({10{received[37]}} & 10'b0101110011) ^ ({10{received[38]}} & 10'b1110001010) ^ ({10{received[39]}} & 10'b0001101111) ^ ({10{received[40]}} & 10'b1101111000) ^ ({10{received[41]}} & 10'b1111110110) ^ ({10{received[42]}} & 10'b1110001111) ^ ({10{received[43]}} & 10'b0001000111) ^ ({10{received[44]}} & 10'b1000111000) ^ ({10{received[45]}} & 10'b0111100100) ^ ({10{received[46]}} & 10'b1100111011) ^ ({10{received[47]}} & 10'b0111101110) ^ ({10{received[48]}} & 10'b1101101011) ^ ({10{received[49]}} & 10'b1101101110) ^ ({10{received[50]}} & 10'b1101000110) ^ ({10{received[51]}} & 10'b1000000110) ^ ({10{received[52]}} & 10'b0000010100) ^ ({10{received[53]}} & 10'b0010100000) ^ ({10{received[54]}} & 10'b0100001001) ^ ({10{received[55]}} & 10'b0001011010) ^ ({10{received[56]}} & 10'b1011010000) ^ ({10{received[57]}} & 10'b1010101101) ^ ({10{received[58]}} & 10'b0101000101) ^ ({10{received[59]}} & 10'b1000111010) ^ ({10{received[60]}} & 10'b0111110100) ^ ({10{received[61]}} & 10'b1110111011) ^ ({10{received[62]}} & 10'b0111100111) ^ ({10{received[63]}} & 10'b1100100011) ^ ({10{received[64]}} & 10'b0100101110) ^ ({10{received[65]}} & 10'b0101100010) ^ ({10{received[66]}} & 10'b1100000010) ^ ({10{received[67]}} & 10'b0000100110) ^ ({10{received[68]}} & 10'b0100110000) ^ ({10{received[69]}} & 10'b0110010010) ^ ({10{received[70]}} & 10'b0010001011) ^ ({10{received[71]}} & 10'b0001010001) ^ ({10{received[72]}} & 10'b1010001000) ^ ({10{received[73]}} & 10'b0001101101) ^ ({10{received[74]}} & 10'b1101101000) ^ ({10{received[75]}} & 10'b1101110110) ^ ({10{received[76]}} & 10'b1110000110) ^ ({10{received[77]}} & 10'b0000001111) ^ ({10{received[78]}} & 10'b0001111000) ^ ({10{received[79]}} & 10'b1111000000) ^ ({10{received[80]}} & 10'b1000111111) ^ ({10{received[81]}} & 10'b0111011100) ^ ({10{received[82]}} & 10'b1011111011) ^ ({10{received[83]}} & 10'b1111110101) ^ ({10{received[84]}} & 10'b1110010111) ^ ({10{received[85]}} & 10'b0010000111) ^ ({10{received[86]}} & 10'b0000110001) ^ ({10{received[87]}} & 10'b0110001000) ^ ({10{received[88]}} & 10'b0001011011) ^ ({10{received[89]}} & 10'b1011011000) ^ ({10{received[90]}} & 10'b1011101101) ^ ({10{received[91]}} & 10'b1101000101) ^ ({10{received[92]}} & 10'b1000011110) ^ ({10{received[93]}} & 10'b0011010100) ^ ({10{received[94]}} & 10'b1010101001) ^ ({10{received[95]}} & 10'b0101100101) ^ ({10{received[96]}} & 10'b1100111010) ^ ({10{received[97]}} & 10'b0111100110) ^ ({10{received[98]}} & 10'b1100101011) ^ ({10{received[99]}} & 10'b0101101110) ^ ({10{received[100]}} & 10'b1101100010) ^ ({10{received[101]}} & 10'b1100100110) ^ ({10{received[102]}} & 10'b0100000110) ^ ({10{received[103]}} & 10'b0000100010) ^ ({10{received[104]}} & 10'b0100010000) ^ ({10{received[105]}} & 10'b0010010010) ^ ({10{received[106]}} & 10'b0010011001) ^ ({10{received[107]}} & 10'b0011000001) ^ ({10{received[108]}} & 10'b1000000001) ^ ({10{received[109]}} & 10'b0000101100) ^ ({10{received[110]}} & 10'b0101100000) ^ ({10{received[111]}} & 10'b1100010010) ^ ({10{received[112]}} & 10'b0010100110) ^ ({10{received[113]}} & 10'b0100111001) ^ ({10{received[114]}} & 10'b0111011010) ^ ({10{received[115]}} & 10'b1011001011) ^ ({10{received[116]}} & 10'b1001110101) ^ ({10{received[117]}} & 10'b1110001100) ^ ({10{received[118]}} & 10'b0001011111) ^ ({10{received[119]}} & 10'b1011111000) ^ ({10{received[120]}} & 10'b1111101101) ^ ({10{received[121]}} & 10'b1101010111) ^ ({10{received[122]}} & 10'b1010001110) ^ ({10{received[123]}} & 10'b0001011101) ^ ({10{received[124]}} & 10'b1011101000) ^ ({10{received[125]}} & 10'b1101101101) ^ ({10{received[126]}} & 10'b1101011110) ^ ({10{received[127]}} & 10'b1011000110) ^ ({10{received[128]}} & 10'b1000011101) ^ ({10{received[129]}} & 10'b0011001100) ^ ({10{received[130]}} & 10'b1001101001) ^ ({10{received[131]}} & 10'b1101101100) ^ ({10{received[132]}} & 10'b1101010110) ^ ({10{received[133]}} & 10'b1010000110) ^ ({10{received[134]}} & 10'b0000011101) ^ ({10{received[135]}} & 10'b0011101000) ^ ({10{received[136]}} & 10'b1101001001) ^ ({10{received[137]}} & 10'b1001111110) ^ ({10{received[138]}} & 10'b1111010100) ^ ({10{received[139]}} & 10'b1010011111) ^ ({10{received[140]}} & 10'b0011010101) ^ ({10{received[141]}} & 10'b1010100001) ^ ({10{received[142]}} & 10'b0100100101) ^ ({10{received[143]}} & 10'b0100111010) ^ ({10{received[144]}} & 10'b0111000010) ^ ({10{received[145]}} & 10'b1000001011) ^ ({10{received[146]}} & 10'b0001111100) ^ ({10{received[147]}} & 10'b1111100000) ^ ({10{received[148]}} & 10'b1100111111) ^ ({10{received[149]}} & 10'b0111001110) ^ ({10{received[150]}} & 10'b1001101011) ^ ({10{received[151]}} & 10'b1101111100) ^ ({10{received[152]}} & 10'b1111010110) ^ ({10{received[153]}} & 10'b1010001111) ^ ({10{received[154]}} & 10'b0001010101) ^ ({10{received[155]}} & 10'b1010101000) ^ ({10{received[156]}} & 10'b0101101101) ^ ({10{received[157]}} & 10'b1101111010) ^ ({10{received[158]}} & 10'b1111100110) ^ ({10{received[159]}} & 10'b1100001111) ^ ({10{received[160]}} & 10'b0001001110) ^ ({10{received[161]}} & 10'b1001110000) ^ ({10{received[162]}} & 10'b1110100100) ^ ({10{received[163]}} & 10'b0100011111) ^ ({10{received[164]}} & 10'b0011101010) ^ ({10{received[165]}} & 10'b1101011001) ^ ({10{received[166]}} & 10'b1011111110) ^ ({10{received[167]}} & 10'b1111011101) ^ ({10{received[168]}} & 10'b1011010111) ^ ({10{received[169]}} & 10'b1010010101) ^ ({10{received[170]}} & 10'b0010000101) ^ ({10{received[171]}} & 10'b0000100001) ^ ({10{received[172]}} & 10'b0100001000) ^ ({10{received[173]}} & 10'b0001010010) ^ ({10{received[174]}} & 10'b1010010000) ^ ({10{received[175]}} & 10'b0010101101) ^ ({10{received[176]}} & 10'b0101100001) ^ ({10{received[177]}} & 10'b1100011010) ^ ({10{received[178]}} & 10'b0011100110) ^ ({10{received[179]}} & 10'b1100111001) ^ ({10{received[180]}} & 10'b0111111110) ^ ({10{received[181]}} & 10'b1111101011) ^ ({10{received[182]}} & 10'b1101100111) ^ ({10{received[183]}} & 10'b1100001110) ^ ({10{received[184]}} & 10'b0001000110) ^ ({10{received[185]}} & 10'b1000110000) ^ ({10{received[186]}} & 10'b0110100100) ^ ({10{received[187]}} & 10'b0100111011) ^ ({10{received[188]}} & 10'b0111001010) ^ ({10{received[189]}} & 10'b1001001011) ^ ({10{received[190]}} & 10'b1001111100) ^ ({10{received[191]}} & 10'b1111000100) ^ ({10{received[192]}} & 10'b1000011111) ^ ({10{received[193]}} & 10'b0011011100) ^ ({10{received[194]}} & 10'b1011101001) ^ ({10{received[195]}} & 10'b1101100101) ^ ({10{received[196]}} & 10'b1100011110) ^ ({10{received[197]}} & 10'b0011000110) ^ ({10{received[198]}} & 10'b1000111001) ^ ({10{received[199]}} & 10'b0111101100) ^ ({10{received[200]}} & 10'b1101111011) ^ ({10{received[201]}} & 10'b1111101110) ^ ({10{received[202]}} & 10'b1101001111) ^ ({10{received[203]}} & 10'b1001001110) ^ ({10{received[204]}} & 10'b1001010100) ^ ({10{received[205]}} & 10'b1010000100) ^ ({10{received[206]}} & 10'b0000001101) ^ ({10{received[207]}} & 10'b0001101000) ^ ({10{received[208]}} & 10'b1101000000) ^ ({10{received[209]}} & 10'b1000110110) ^ ({10{received[210]}} & 10'b0110010100) ^ ({10{received[211]}} & 10'b0010111011) ^ ({10{received[212]}} & 10'b0111010001) ^ ({10{received[213]}} & 10'b1010010011) ^ ({10{received[214]}} & 10'b0010110101) ^ ({10{received[215]}} & 10'b0110100001) ^ ({10{received[216]}} & 10'b0100010011) ^ ({10{received[217]}} & 10'b0010001010) ^ ({10{received[218]}} & 10'b0001011001) ^ ({10{received[219]}} & 10'b1011001000) ^ ({10{received[220]}} & 10'b1001101101) ^ ({10{received[221]}} & 10'b1101001100) ^ ({10{received[222]}} & 10'b1001010110) ^ ({10{received[223]}} & 10'b1010010100) ^ ({10{received[224]}} & 10'b0010001101) ^ ({10{received[225]}} & 10'b0001100001) ^ ({10{received[226]}} & 10'b1100001000) ^ ({10{received[227]}} & 10'b0001110110) ^ ({10{received[228]}} & 10'b1110110000) ^ ({10{received[229]}} & 10'b0110111111) ^ ({10{received[230]}} & 10'b0111100011) ^ ({10{received[231]}} & 10'b1100000011) ^ ({10{received[232]}} & 10'b0000101110) ^ ({10{received[233]}} & 10'b0101110000) ^ ({10{received[234]}} & 10'b1110010010) ^ ({10{received[235]}} & 10'b0010101111) ^ ({10{received[236]}} & 10'b0101110001) ^ ({10{received[237]}} & 10'b1110011010) ^ ({10{received[238]}} & 10'b0011101111) ^ ({10{received[239]}} & 10'b1101110001) ^ ({10{received[240]}} & 10'b1110111110) ^ ({10{received[241]}} & 10'b0111001111) ^ ({10{received[242]}} & 10'b1001100011) ^ ({10{received[243]}} & 10'b1100111100) ^ ({10{received[244]}} & 10'b0111010110) ^ ({10{received[245]}} & 10'b1010101011) ^ ({10{received[246]}} & 10'b0101110101) ^ ({10{received[247]}} & 10'b1110111010) ^ ({10{received[248]}} & 10'b0111101111) ^ ({10{received[249]}} & 10'b1101100011) ^ ({10{received[250]}} & 10'b1100101110) ^ ({10{received[251]}} & 10'b0101000110) ^ ({10{received[252]}} & 10'b1000100010) ^ ({10{received[253]}} & 10'b0100110100) ^ ({10{received[254]}} & 10'b0110110010) ^ ({10{received[255]}} & 10'b0110001011) ^ ({10{received[256]}} & 10'b0001000011) ^ ({10{received[257]}} & 10'b1000011000) ^ ({10{received[258]}} & 10'b0011100100) ^ ({10{received[259]}} & 10'b1100101001) ^ ({10{received[260]}} & 10'b0101111110) ^ ({10{received[261]}} & 10'b1111100010) ^ ({10{received[262]}} & 10'b1100101111) ^ ({10{received[263]}} & 10'b0101001110) ^ ({10{received[264]}} & 10'b1001100010) ^ ({10{received[265]}} & 10'b1100110100) ^ ({10{received[266]}} & 10'b0110010110) ^ ({10{received[267]}} & 10'b0010101011) ^ ({10{received[268]}} & 10'b0101010001) ^ ({10{received[269]}} & 10'b1010011010) ^ ({10{received[270]}} & 10'b0011111101) ^ ({10{received[271]}} & 10'b1111100001) ^ ({10{received[272]}} & 10'b1100110111) ^ ({10{received[273]}} & 10'b0110001110) ^ ({10{received[274]}} & 10'b0001101011) ^ ({10{received[275]}} & 10'b1101011000) ^ ({10{received[276]}} & 10'b1011110110) ^ ({10{received[277]}} & 10'b1110011101) ^ ({10{received[278]}} & 10'b0011010111) ^ ({10{received[279]}} & 10'b1010110001) ^ ({10{received[280]}} & 10'b0110100101) ^ ({10{received[281]}} & 10'b0100110011) ^ ({10{received[282]}} & 10'b0110001010) ^ ({10{received[283]}} & 10'b0001001011) ^ ({10{received[284]}} & 10'b1001011000) ^ ({10{received[285]}} & 10'b1011100100) ^ ({10{received[286]}} & 10'b1100001101) ^ ({10{received[287]}} & 10'b0001011110) ^ ({10{received[288]}} & 10'b1011110000) ^ ({10{received[289]}} & 10'b1110101101) ^ ({10{received[290]}} & 10'b0101010111) ^ ({10{received[291]}} & 10'b1010101010) ^ ({10{received[292]}} & 10'b0101111101) ^ ({10{received[293]}} & 10'b1111111010) ^ ({10{received[294]}} & 10'b1111101111) ^ ({10{received[295]}} & 10'b1101000111) ^ ({10{received[296]}} & 10'b1000001110) ^ ({10{received[297]}} & 10'b0001010100) ^ ({10{received[298]}} & 10'b1010100000) ^ ({10{received[299]}} & 10'b0100101101) ^ ({10{received[300]}} & 10'b0101111010) ^ ({10{received[301]}} & 10'b1111000010) ^ ({10{received[302]}} & 10'b1000101111) ^ ({10{received[303]}} & 10'b0101011100) ^ ({10{received[304]}} & 10'b1011110010) ^ ({10{received[305]}} & 10'b1110111101) ^ ({10{received[306]}} & 10'b0111010111) ^ ({10{received[307]}} & 10'b1010100011) ^ ({10{received[308]}} & 10'b0100110101) ^ ({10{received[309]}} & 10'b0110111010) ^ ({10{received[310]}} & 10'b0111001011) ^ ({10{received[311]}} & 10'b1001000011) ^ ({10{received[312]}} & 10'b1000111100) ^ ({10{received[313]}} & 10'b0111000100) ^ ({10{received[314]}} & 10'b1000111011) ^ ({10{received[315]}} & 10'b0111111100) ^ ({10{received[316]}} & 10'b1111111011) ^ ({10{received[317]}} & 10'b1111100111) ^ ({10{received[318]}} & 10'b1100000111) ^ ({10{received[319]}} & 10'b0000001110) ^ ({10{received[320]}} & 10'b0001110000) ^ ({10{received[321]}} & 10'b1110000000) ^ ({10{received[322]}} & 10'b0000111111) ^ ({10{received[323]}} & 10'b0111111000) ^ ({10{received[324]}} & 10'b1111011011) ^ ({10{received[325]}} & 10'b1011100111) ^ ({10{received[326]}} & 10'b1100010101) ^ ({10{received[327]}} & 10'b0010011110) ^ ({10{received[328]}} & 10'b0011111001) ^ ({10{received[329]}} & 10'b1111000001) ^ ({10{received[330]}} & 10'b1000110111) ^ ({10{received[331]}} & 10'b0110011100) ^ ({10{received[332]}} & 10'b0011111011) ^ ({10{received[333]}} & 10'b1111010001) ^ ({10{received[334]}} & 10'b1010110111) ^ ({10{received[335]}} & 10'b0110010101) ^ ({10{received[336]}} & 10'b0010110011) ^ ({10{received[337]}} & 10'b0110010001) ^ ({10{received[338]}} & 10'b0010010011) ^ ({10{received[339]}} & 10'b0010010001) ^ ({10{received[340]}} & 10'b0010000001) ^ ({10{received[341]}} & 10'b0000000001) ^ ({10{received[342]}} & 10'b0000001000) ^ ({10{received[343]}} & 10'b0001000000) ^ ({10{received[344]}} & 10'b1000000000) ^ ({10{received[345]}} & 10'b0000100100) ^ ({10{received[346]}} & 10'b0100100000) ^ ({10{received[347]}} & 10'b0100010010) ^ ({10{received[348]}} & 10'b0010000010) ^ ({10{received[349]}} & 10'b0000011001) ^ ({10{received[350]}} & 10'b0011001000) ^ ({10{received[351]}} & 10'b1001001001) ^ ({10{received[352]}} & 10'b1001101100) ^ ({10{received[353]}} & 10'b1101000100) ^ ({10{received[354]}} & 10'b1000010110) ^ ({10{received[355]}} & 10'b0010010100) ^ ({10{received[356]}} & 10'b0010101001) ^ ({10{received[357]}} & 10'b0101000001) ^ ({10{received[358]}} & 10'b1000011010) ^ ({10{received[359]}} & 10'b0011110100) ^ ({10{received[360]}} & 10'b1110101001) ^ ({10{received[361]}} & 10'b0101110111) ^ ({10{received[362]}} & 10'b1110101010) ^ ({10{received[363]}} & 10'b0101101111) ^ ({10{received[364]}} & 10'b1101101010) ^ ({10{received[365]}} & 10'b1101100110) ^ ({10{received[366]}} & 10'b1100000110) ^ ({10{received[367]}} & 10'b0000000110) ^ ({10{received[368]}} & 10'b0000110000) ^ ({10{received[369]}} & 10'b0110000000) ^ ({10{received[370]}} & 10'b0000011011) ^ ({10{received[371]}} & 10'b0011011000) ^ ({10{received[372]}} & 10'b1011001001) ^ ({10{received[373]}} & 10'b1001100101) ^ ({10{received[374]}} & 10'b1100001100) ^ ({10{received[375]}} & 10'b0001010110) ^ ({10{received[376]}} & 10'b1010110000) ^ ({10{received[377]}} & 10'b0110101101) ^ ({10{received[378]}} & 10'b0101110011) ^ ({10{received[379]}} & 10'b1110001010) ^ ({10{received[380]}} & 10'b0001101111) ^ ({10{received[381]}} & 10'b1101111000) ^ ({10{received[382]}} & 10'b1111110110) ^ ({10{received[383]}} & 10'b1110001111) ^ ({10{received[384]}} & 10'b0001000111) ^ ({10{received[385]}} & 10'b1000111000) ^ ({10{received[386]}} & 10'b0111100100) ^ ({10{received[387]}} & 10'b1100111011) ^ ({10{received[388]}} & 10'b0111101110) ^ ({10{received[389]}} & 10'b1101101011) ^ ({10{received[390]}} & 10'b1101101110) ^ ({10{received[391]}} & 10'b1101000110) ^ ({10{received[392]}} & 10'b1000000110) ^ ({10{received[393]}} & 10'b0000010100) ^ ({10{received[394]}} & 10'b0010100000) ^ ({10{received[395]}} & 10'b0100001001) ^ ({10{received[396]}} & 10'b0001011010) ^ ({10{received[397]}} & 10'b1011010000) ^ ({10{received[398]}} & 10'b1010101101) ^ ({10{received[399]}} & 10'b0101000101) ^ ({10{received[400]}} & 10'b1000111010) ^ ({10{received[401]}} & 10'b0111110100) ^ ({10{received[402]}} & 10'b1110111011) ^ ({10{received[403]}} & 10'b0111100111) ^ ({10{received[404]}} & 10'b1100100011) ^ ({10{received[405]}} & 10'b0100101110) ^ ({10{received[406]}} & 10'b0101100010) ^ ({10{received[407]}} & 10'b1100000010) ^ ({10{received[408]}} & 10'b0000100110) ^ ({10{received[409]}} & 10'b0100110000) ^ ({10{received[410]}} & 10'b0110010010) ^ ({10{received[411]}} & 10'b0010001011) ^ ({10{received[412]}} & 10'b0001010001) ^ ({10{received[413]}} & 10'b1010001000) ^ ({10{received[414]}} & 10'b0001101101) ^ ({10{received[415]}} & 10'b1101101000) ^ ({10{received[416]}} & 10'b1101110110) ^ ({10{received[417]}} & 10'b1110000110) ^ ({10{received[418]}} & 10'b0000001111) ^ ({10{received[419]}} & 10'b0001111000) ^ ({10{received[420]}} & 10'b1111000000) ^ ({10{received[421]}} & 10'b1000111111) ^ ({10{received[422]}} & 10'b0111011100) ^ ({10{received[423]}} & 10'b1011111011) ^ ({10{received[424]}} & 10'b1111110101) ^ ({10{received[425]}} & 10'b1110010111) ^ ({10{received[426]}} & 10'b0010000111) ^ ({10{received[427]}} & 10'b0000110001) ^ ({10{received[428]}} & 10'b0110001000) ^ ({10{received[429]}} & 10'b0001011011) ^ ({10{received[430]}} & 10'b1011011000) ^ ({10{received[431]}} & 10'b1011101101) ^ ({10{received[432]}} & 10'b1101000101) ^ ({10{received[433]}} & 10'b1000011110) ^ ({10{received[434]}} & 10'b0011010100) ^ ({10{received[435]}} & 10'b1010101001) ^ ({10{received[436]}} & 10'b0101100101) ^ ({10{received[437]}} & 10'b1100111010) ^ ({10{received[438]}} & 10'b0111100110) ^ ({10{received[439]}} & 10'b1100101011) ^ ({10{received[440]}} & 10'b0101101110) ^ ({10{received[441]}} & 10'b1101100010) ^ ({10{received[442]}} & 10'b1100100110) ^ ({10{received[443]}} & 10'b0100000110) ^ ({10{received[444]}} & 10'b0000100010) ^ ({10{received[445]}} & 10'b0100010000) ^ ({10{received[446]}} & 10'b0010010010) ^ ({10{received[447]}} & 10'b0010011001) ^ ({10{received[448]}} & 10'b0011000001) ^ ({10{received[449]}} & 10'b1000000001) ^ ({10{received[450]}} & 10'b0000101100) ^ ({10{received[451]}} & 10'b0101100000) ^ ({10{received[452]}} & 10'b1100010010) ^ ({10{received[453]}} & 10'b0010100110) ^ ({10{received[454]}} & 10'b0100111001) ^ ({10{received[455]}} & 10'b0111011010) ^ ({10{received[456]}} & 10'b1011001011) ^ ({10{received[457]}} & 10'b1001110101) ^ ({10{received[458]}} & 10'b1110001100) ^ ({10{received[459]}} & 10'b0001011111) ^ ({10{received[460]}} & 10'b1011111000) ^ ({10{received[461]}} & 10'b1111101101) ^ ({10{received[462]}} & 10'b1101010111) ^ ({10{received[463]}} & 10'b1010001110) ^ ({10{received[464]}} & 10'b0001011101) ^ ({10{received[465]}} & 10'b1011101000) ^ ({10{received[466]}} & 10'b1101101101) ^ ({10{received[467]}} & 10'b1101011110) ^ ({10{received[468]}} & 10'b1011000110) ^ ({10{received[469]}} & 10'b1000011101) ^ ({10{received[470]}} & 10'b0011001100) ^ ({10{received[471]}} & 10'b1001101001) ^ ({10{received[472]}} & 10'b1101101100) ^ ({10{received[473]}} & 10'b1101010110) ^ ({10{received[474]}} & 10'b1010000110) ^ ({10{received[475]}} & 10'b0000011101) ^ ({10{received[476]}} & 10'b0011101000) ^ ({10{received[477]}} & 10'b1101001001) ^ ({10{received[478]}} & 10'b1001111110) ^ ({10{received[479]}} & 10'b1111010100) ^ ({10{received[480]}} & 10'b1010011111) ^ ({10{received[481]}} & 10'b0011010101) ^ ({10{received[482]}} & 10'b1010100001) ^ ({10{received[483]}} & 10'b0100100101) ^ ({10{received[484]}} & 10'b0100111010) ^ ({10{received[485]}} & 10'b0111000010) ^ ({10{received[486]}} & 10'b1000001011) ^ ({10{received[487]}} & 10'b0001111100) ^ ({10{received[488]}} & 10'b1111100000) ^ ({10{received[489]}} & 10'b1100111111) ^ ({10{received[490]}} & 10'b0111001110) ^ ({10{received[491]}} & 10'b1001101011) ^ ({10{received[492]}} & 10'b1101111100) ^ ({10{received[493]}} & 10'b1111010110) ^ ({10{received[494]}} & 10'b1010001111) ^ ({10{received[495]}} & 10'b0001010101) ^ ({10{received[496]}} & 10'b1010101000) ^ ({10{received[497]}} & 10'b0101101101) ^ ({10{received[498]}} & 10'b1101111010) ^ ({10{received[499]}} & 10'b1111100110) ^ ({10{received[500]}} & 10'b1100001111) ^ ({10{received[501]}} & 10'b0001001110) ^ ({10{received[502]}} & 10'b1001110000) ^ ({10{received[503]}} & 10'b1110100100) ^ ({10{received[504]}} & 10'b0100011111) ^ ({10{received[505]}} & 10'b0011101010) ^ ({10{received[506]}} & 10'b1101011001) ^ ({10{received[507]}} & 10'b1011111110) ^ ({10{received[508]}} & 10'b1111011101) ^ ({10{received[509]}} & 10'b1011010111) ^ ({10{received[510]}} & 10'b1010010101) ^ ({10{received[511]}} & 10'b0010000101) ^ ({10{received[512]}} & 10'b0000100001) ^ ({10{received[513]}} & 10'b0100001000) ^ ({10{received[514]}} & 10'b0001010010) ^ ({10{received[515]}} & 10'b1010010000) ^ ({10{received[516]}} & 10'b0010101101) ^ ({10{received[517]}} & 10'b0101100001) ^ ({10{received[518]}} & 10'b1100011010) ^ ({10{received[519]}} & 10'b0011100110) ^ ({10{received[520]}} & 10'b1100111001) ^ ({10{received[521]}} & 10'b0111111110) ^ ({10{received[522]}} & 10'b1111101011) ^ ({10{received[523]}} & 10'b1101100111) ^ ({10{received[524]}} & 10'b1100001110) ^ ({10{received[525]}} & 10'b0001000110) ^ ({10{received[526]}} & 10'b1000110000) ^ ({10{received[527]}} & 10'b0110100100) ^ ({10{received[528]}} & 10'b0100111011) ^ ({10{received[529]}} & 10'b0111001010) ^ ({10{received[530]}} & 10'b1001001011) ^ ({10{received[531]}} & 10'b1001111100) ^ ({10{received[532]}} & 10'b1111000100) ^ ({10{received[533]}} & 10'b1000011111) ^ ({10{received[534]}} & 10'b0011011100) ^ ({10{received[535]}} & 10'b1011101001) ^ ({10{received[536]}} & 10'b1101100101) ^ ({10{received[537]}} & 10'b1100011110) ^ ({10{received[538]}} & 10'b0011000110) ^ ({10{received[539]}} & 10'b1000111001) ^ ({10{received[540]}} & 10'b0111101100) ^ ({10{received[541]}} & 10'b1101111011);
  assign syndrome4 = ({10{received[0]}} & 10'b0000000001) ^ 
  ({10{received[1]}} & 10'b0000010000) ^ ({10{received[2]}} & 10'b0100000000) ^ ({10{received[3]}} & 10'b0000100100) ^ ({10{received[4]}} & 10'b1001000000) ^ ({10{received[5]}} & 10'b0001000001) ^ ({10{received[6]}} & 10'b0000011001) ^ ({10{received[7]}} & 10'b0110010000) ^ ({10{received[8]}} & 10'b0100110110) ^ ({10{received[9]}} & 10'b1101000100) ^ ({10{received[10]}} & 10'b0000100101) ^ ({10{received[11]}} & 10'b1001010000) ^ ({10{received[12]}} & 10'b0101000001) ^ ({10{received[13]}} & 10'b0000111101) ^ ({10{received[14]}} & 10'b1111010000) ^ ({10{received[15]}} & 10'b0101110111) ^ ({10{received[16]}} & 10'b1101011101) ^ ({10{received[17]}} & 10'b0110110101) ^ ({10{received[18]}} & 10'b1101100110) ^ ({10{received[19]}} & 10'b1000000101) ^ ({10{received[20]}} & 10'b0000011000) ^ ({10{received[21]}} & 10'b0110000000) ^ ({10{received[22]}} & 10'b0000110110) ^ ({10{received[23]}} & 10'b1101100000) ^ ({10{received[24]}} & 10'b1001100101) ^ ({10{received[25]}} & 10'b1000010001) ^ ({10{received[26]}} & 10'b0101011000) ^ ({10{received[27]}} & 10'b0110101101) ^ ({10{received[28]}} & 10'b1011100110) ^ ({10{received[29]}} & 10'b1000110011) ^ ({10{received[30]}} & 10'b1101111000) ^ ({10{received[31]}} & 10'b1111100101) ^ ({10{received[32]}} & 10'b1000100111) ^ ({10{received[33]}} & 10'b1000111000) ^ ({10{received[34]}} & 10'b1111001000) ^ ({10{received[35]}} & 10'b0011110111) ^ ({10{received[36]}} & 10'b1101101011) ^ ({10{received[37]}} & 10'b1011010101) ^ ({10{received[38]}} & 10'b0100000011) ^ ({10{received[39]}} & 10'b0000010100) ^ ({10{received[40]}} & 10'b0101000000) ^ ({10{received[41]}} & 10'b0000101101) ^ ({10{received[42]}} & 10'b1011010000) ^ ({10{received[43]}} & 10'b0101010011) ^ ({10{received[44]}} & 10'b0100011101) ^ ({10{received[45]}} & 10'b0111110100) ^ ({10{received[46]}} & 10'b1101111111) ^ ({10{received[47]}} & 10'b1110010101) ^ ({10{received[48]}} & 10'b0100101110) ^ ({10{received[49]}} & 10'b1011000100) ^ ({10{received[50]}} & 10'b0000010011) ^ ({10{received[51]}} & 10'b0100110000) ^ ({10{received[52]}} & 10'b1100100100) ^ ({10{received[53]}} & 10'b1000101100) ^ ({10{received[54]}} & 10'b1010001000) ^ ({10{received[55]}} & 10'b0011011010) ^ ({10{received[56]}} & 10'b0110111011) ^ ({10{received[57]}} & 10'b1110000110) ^ ({10{received[58]}} & 10'b0000011110) ^ ({10{received[59]}} & 10'b0111100000) ^ ({10{received[60]}} & 10'b1000111111) ^ ({10{received[61]}} & 10'b1110111000) ^ ({10{received[62]}} & 10'b1111111110) ^ ({10{received[63]}} & 10'b1110010111) ^ ({10{received[64]}} & 10'b0100001110) ^ ({10{received[65]}} & 10'b0011000100) ^ ({10{received[66]}} & 10'b0001011011) ^ ({10{received[67]}} & 10'b0110111001) ^ ({10{received[68]}} & 10'b1110100110) ^ ({10{received[69]}} & 10'b1000011110) ^ ({10{received[70]}} & 10'b0110101000) ^ ({10{received[71]}} & 10'b1010110110) ^ ({10{received[72]}} & 10'b1100111010) ^ ({10{received[73]}} & 10'b1111001100) ^ ({10{received[74]}} & 10'b0010110111) ^ ({10{received[75]}} & 10'b1101100010) ^ ({10{received[76]}} & 10'b1001000101) ^ ({10{received[77]}} & 10'b0000010001) ^ ({10{received[78]}} & 10'b0100010000) ^ ({10{received[79]}} & 10'b0100100100) ^ ({10{received[80]}} & 10'b1001100100) ^ ({10{received[81]}} & 10'b1000000001) ^ ({10{received[82]}} & 10'b0001011000) ^ ({10{received[83]}} & 10'b0110001001) ^ ({10{received[84]}} & 10'b0010100110) ^ ({10{received[85]}} & 10'b1001110010) ^ ({10{received[86]}} & 10'b1101100001) ^ ({10{received[87]}} & 10'b1001110101) ^ ({10{received[88]}} & 10'b1100010001) ^ ({10{received[89]}} & 10'b0101111100) ^ ({10{received[90]}} & 10'b1111101101) ^ ({10{received[91]}} & 10'b1010100111) ^ ({10{received[92]}} & 10'b1000101010) ^ ({10{received[93]}} & 10'b1011101000) ^ ({10{received[94]}} & 10'b1011010011) ^ ({10{received[95]}} & 10'b0101100011) ^ ({10{received[96]}} & 10'b1000011101) ^ ({10{received[97]}} & 10'b0110011000) ^ ({10{received[98]}} & 10'b0110110110) ^ ({10{received[99]}} & 10'b1101010110) ^ ({10{received[100]}} & 10'b0100000101) ^ ({10{received[101]}} & 10'b0001110100) ^ ({10{received[102]}} & 10'b1101001001) ^ ({10{received[103]}} & 10'b0011110101) ^ ({10{received[104]}} & 10'b1101001011) ^ ({10{received[105]}} & 10'b0011010101) ^ ({10{received[106]}} & 10'b0101001011) ^ ({10{received[107]}} & 10'b0010011101) ^ ({10{received[108]}} & 10'b0111000010) ^ ({10{received[109]}} & 10'b0000011111) ^ ({10{received[110]}} & 10'b0111110000) ^ ({10{received[111]}} & 10'b1100111111) ^ ({10{received[112]}} & 10'b1110011100) ^ ({10{received[113]}} & 10'b0110111110) ^ ({10{received[114]}} & 10'b1111010110) ^ ({10{received[115]}} & 10'b0100010111) ^ ({10{received[116]}} & 10'b0101010100) ^ ({10{received[117]}} & 10'b0101101101) ^ ({10{received[118]}} & 10'b1011111101) ^ ({10{received[119]}} & 10'b1110000011) ^ ({10{received[120]}} & 10'b0001001110) ^ ({10{received[121]}} & 10'b0011101001) ^ ({10{received[122]}} & 10'b1010001011) ^ ({10{received[123]}} & 10'b0011101010) ^ ({10{received[124]}} & 10'b1010111011) ^ ({10{received[125]}} & 10'b1111101010) ^ ({10{received[126]}} & 10'b1011010111) ^ ({10{received[127]}} & 10'b0100100011) ^ ({10{received[128]}} & 10'b1000010100) ^ ({10{received[129]}} & 10'b0100001000) ^ ({10{received[130]}} & 10'b0010100100) ^ ({10{received[131]}} & 10'b1001010010) ^ ({10{received[132]}} & 10'b0101100001) ^ ({10{received[133]}} & 10'b1000111101) ^ ({10{received[134]}} & 10'b1110011000) ^ ({10{received[135]}} & 10'b0111111110) ^ ({10{received[136]}} & 10'b1111011111) ^ ({10{received[137]}} & 10'b0110000111) ^ ({10{received[138]}} & 10'b0001000110) ^ ({10{received[139]}} & 10'b0001101001) ^ ({10{received[140]}} & 10'b1010011001) ^ ({10{received[141]}} & 10'b0111001010) ^ ({10{received[142]}} & 10'b0010011111) ^ ({10{received[143]}} & 10'b0111100010) ^ ({10{received[144]}} & 10'b1000011111) ^ ({10{received[145]}} & 10'b0110111000) ^ ({10{received[146]}} & 10'b1110110110) ^ ({10{received[147]}} & 10'b1100011110) ^ ({10{received[148]}} & 10'b0110001100) ^ ({10{received[149]}} & 10'b0011110110) ^ ({10{received[150]}} & 10'b1101111011) ^ ({10{received[151]}} & 10'b1111010101) ^ ({10{received[152]}} & 10'b0100100111) ^ ({10{received[153]}} & 10'b1001010100) ^ ({10{received[154]}} & 10'b0100000001) ^ ({10{received[155]}} & 10'b0000110100) ^ ({10{received[156]}} & 10'b1101000000) ^ ({10{received[157]}} & 10'b0001100101) ^ ({10{received[158]}} & 10'b1001011001) ^ ({10{received[159]}} & 10'b0111010001) ^ ({10{received[160]}} & 10'b0100101111) ^ ({10{received[161]}} & 10'b1011010100) ^ ({10{received[162]}} & 10'b0100010011) ^ ({10{received[163]}} & 10'b0100010100) ^ ({10{received[164]}} & 10'b0101100100) ^ ({10{received[165]}} & 10'b1001101101) ^ ({10{received[166]}} & 10'b1010010001) ^ ({10{received[167]}} & 10'b0101001010) ^ ({10{received[168]}} & 10'b0010001101) ^ ({10{received[169]}} & 10'b0011000010) ^ ({10{received[170]}} & 10'b0000111011) ^ ({10{received[171]}} & 10'b1110110000) ^ ({10{received[172]}} & 10'b1101111110) ^ ({10{received[173]}} & 10'b1110000101) ^ ({10{received[174]}} & 10'b0000101110) ^ ({10{received[175]}} & 10'b1011100000) ^ ({10{received[176]}} & 10'b1001010011) ^ ({10{received[177]}} & 10'b0101110001) ^ ({10{received[178]}} & 10'b1100111101) ^ ({10{received[179]}} & 10'b1110111100) ^ ({10{received[180]}} & 10'b1110111110) ^ ({10{received[181]}} & 10'b1110011110) ^ ({10{received[182]}} & 10'b0110011110) ^ ({10{received[183]}} & 10'b0111010110) ^ ({10{received[184]}} & 10'b0101011111) ^ ({10{received[185]}} & 10'b0111011101) ^ ({10{received[186]}} & 10'b0111101111) ^ ({10{received[187]}} & 10'b1011001111) ^ ({10{received[188]}} & 10'b0010100011) ^ ({10{received[189]}} & 10'b1000100010) ^ ({10{received[190]}} & 10'b1001101000) ^ ({10{received[191]}} & 10'b1011000001) ^ ({10{received[192]}} & 10'b0001000011) ^ ({10{received[193]}} & 10'b0000111001) ^ ({10{received[194]}} & 10'b1110010000) ^ ({10{received[195]}} & 10'b0101111110) ^ ({10{received[196]}} & 10'b1111001101) ^ ({10{received[197]}} & 10'b0010100111) ^ ({10{received[198]}} & 10'b1001100010) ^ ({10{received[199]}} & 10'b1001100001) ^ ({10{received[200]}} & 10'b1001010001) ^ ({10{received[201]}} & 10'b0101010001) ^ ({10{received[202]}} & 10'b0100111101) ^ ({10{received[203]}} & 10'b1111110100) ^ ({10{received[204]}} & 10'b1100110111) ^ ({10{received[205]}} & 10'b1100011100) ^ ({10{received[206]}} & 10'b0110101100) ^ ({10{received[207]}} & 10'b1011110110) ^ ({10{received[208]}} & 10'b1100110011) ^ ({10{received[209]}} & 10'b1101011100) ^ ({10{received[210]}} & 10'b0110100101) ^ ({10{received[211]}} & 10'b1001100110) ^ ({10{received[212]}} & 10'b1000100001) ^ ({10{received[213]}} & 10'b1001011000) ^ ({10{received[214]}} & 10'b0111000001) ^ ({10{received[215]}} & 10'b0000101111) ^ ({10{received[216]}} & 10'b1011110000) ^ ({10{received[217]}} & 10'b1101010011) ^ ({10{received[218]}} & 10'b0101010101) ^ ({10{received[219]}} & 10'b0101111101) ^ ({10{received[220]}} & 10'b1111111101) ^ ({10{received[221]}} & 10'b1110100111) ^ ({10{received[222]}} & 10'b1000001110) ^ ({10{received[223]}} & 10'b0010101000) ^ ({10{received[224]}} & 10'b1010010010) ^ ({10{received[225]}} & 10'b0101111010) ^ ({10{received[226]}} & 10'b1110001101) ^ ({10{received[227]}} & 10'b0010101110) ^ ({10{received[228]}} & 10'b1011110010) ^ ({10{received[229]}} & 10'b1101110011) ^ ({10{received[230]}} & 10'b1101010101) ^ ({10{received[231]}} & 10'b0100110101) ^ ({10{received[232]}} & 10'b1101110100) ^ ({10{received[233]}} & 10'b1100100101) ^ ({10{received[234]}} & 10'b1000111100) ^ ({10{received[235]}} & 10'b1110001000) ^ ({10{received[236]}} & 10'b0011111110) ^ ({10{received[237]}} & 10'b1111111011) ^ ({10{received[238]}} & 10'b1111000111) ^ ({10{received[239]}} & 10'b0000000111) ^ ({10{received[240]}} & 10'b0001110000) ^ ({10{received[241]}} & 10'b1100001001) ^ ({10{received[242]}} & 10'b0011111100) ^ ({10{received[243]}} & 10'b1111011011) ^ ({10{received[244]}} & 10'b0111000111) ^ ({10{received[245]}} & 10'b0001001111) ^ ({10{received[246]}} & 10'b0011111001) ^ ({10{received[247]}} & 10'b1110001011) ^ ({10{received[248]}} & 10'b0011001110) ^ ({10{received[249]}} & 10'b0011111011) ^ ({10{received[250]}} & 10'b1110101011) ^ ({10{received[251]}} & 10'b1011001110) ^ ({10{received[252]}} & 10'b0010110011) ^ ({10{received[253]}} & 10'b1100100010) ^ ({10{received[254]}} & 10'b1001001100) ^ ({10{received[255]}} & 10'b0010000001) ^ ({10{received[256]}} & 10'b0000000010) ^ ({10{received[257]}} & 10'b0000100000) ^ ({10{received[258]}} & 10'b1000000000) ^ ({10{received[259]}} & 10'b0001001000) ^ ({10{received[260]}} & 10'b0010001001) ^ ({10{received[261]}} & 10'b0010000010) ^ ({10{received[262]}} & 10'b0000110010) ^ ({10{received[263]}} & 10'b1100100000) ^ ({10{received[264]}} & 10'b1001101100) ^ ({10{received[265]}} & 10'b1010000001) ^ ({10{received[266]}} & 10'b0001001010) ^ ({10{received[267]}} & 10'b0010101001) ^ ({10{received[268]}} & 10'b1010000010) ^ ({10{received[269]}} & 10'b0001111010) ^ ({10{received[270]}} & 10'b1110101001) ^ ({10{received[271]}} & 10'b1011101110) ^ ({10{received[272]}} & 10'b1010110011) ^ ({10{received[273]}} & 10'b1101101010) ^ ({10{received[274]}} & 10'b1011000101) ^ ({10{received[275]}} & 10'b0000000011) ^ ({10{received[276]}} & 10'b0000110000) ^ ({10{received[277]}} & 10'b1100000000) ^ ({10{received[278]}} & 10'b0001101100) ^ ({10{received[279]}} & 10'b1011001001) ^ ({10{received[280]}} & 10'b0011000011) ^ ({10{received[281]}} & 10'b0000101011) ^ ({10{received[282]}} & 10'b1010110000) ^ ({10{received[283]}} & 10'b1101011010) ^ ({10{received[284]}} & 10'b0111000101) ^ ({10{received[285]}} & 10'b0001101111) ^ ({10{received[286]}} & 10'b1011111001) ^ ({10{received[287]}} & 10'b1111000011) ^ ({10{received[288]}} & 10'b0001000111) ^ ({10{received[289]}} & 10'b0001111001) ^ ({10{received[290]}} & 10'b1110011001) ^ ({10{received[291]}} & 10'b0111101110) ^ ({10{received[292]}} & 10'b1011011111) ^ ({10{received[293]}} & 10'b0110100011) ^ ({10{received[294]}} & 10'b1000000110) ^ ({10{received[295]}} & 10'b0000101000) ^ ({10{received[296]}} & 10'b1010000000) ^ ({10{received[297]}} & 10'b0001011010) ^ ({10{received[298]}} & 10'b0110101001) ^ ({10{received[299]}} & 10'b1010100110) ^ ({10{received[300]}} & 10'b1000111010) ^ ({10{received[301]}} & 10'b1111101000) ^ ({10{received[302]}} & 10'b1011110111) ^ ({10{received[303]}} & 10'b1100100011) ^ ({10{received[304]}} & 10'b1001011100) ^ ({10{received[305]}} & 10'b0110000001) ^ ({10{received[306]}} & 10'b0000100110) ^ ({10{received[307]}} & 10'b1001100000) ^ ({10{received[308]}} & 10'b1001000001) ^ ({10{received[309]}} & 10'b0001010001) ^ ({10{received[310]}} & 10'b0100011001) ^ ({10{received[311]}} & 10'b0110110100) ^ ({10{received[312]}} & 10'b1101110110) ^ ({10{received[313]}} & 10'b1100000101) ^ ({10{received[314]}} & 10'b0000111100) ^ ({10{received[315]}} & 10'b1111000000) ^ ({10{received[316]}} & 10'b0001110111) ^ ({10{received[317]}} & 10'b1101111001) ^ ({10{received[318]}} & 10'b1111110101) ^ ({10{received[319]}} & 10'b1100100111) ^ ({10{received[320]}} & 10'b1000011100) ^ ({10{received[321]}} & 10'b0110001000) ^ ({10{received[322]}} & 10'b0010110110) ^ ({10{received[323]}} & 10'b1101110010) ^ ({10{received[324]}} & 10'b1101000101) ^ ({10{received[325]}} & 10'b0000110101) ^ ({10{received[326]}} & 10'b1101010000) ^ ({10{received[327]}} & 10'b0101100101) ^ ({10{received[328]}} & 10'b1001111101) ^ ({10{received[329]}} & 10'b1110010001) ^ ({10{received[330]}} & 10'b0101101110) ^ ({10{received[331]}} & 10'b1011001101) ^ ({10{received[332]}} & 10'b0010000011) ^ ({10{received[333]}} & 10'b0000100010) ^ ({10{received[334]}} & 10'b1000100000) ^ ({10{received[335]}} & 10'b1001001000) ^ ({10{received[336]}} & 10'b0011000001) ^ ({10{received[337]}} & 10'b0000001011) ^ ({10{received[338]}} & 10'b0010110000) ^ ({10{received[339]}} & 10'b1100010010) ^ ({10{received[340]}} & 10'b0101001100) ^ ({10{received[341]}} & 10'b0011101101) ^ ({10{received[342]}} & 10'b1011001011) ^ ({10{received[343]}} & 10'b0011100011) ^ ({10{received[344]}} & 10'b1000101011) ^ ({10{received[345]}} & 10'b1011111000) ^ ({10{received[346]}} & 10'b1111010011) ^ ({10{received[347]}} & 10'b0101000111) ^ ({10{received[348]}} & 10'b0001011101) ^ ({10{received[349]}} & 10'b0111011001) ^ ({10{received[350]}} & 10'b0110101111) ^ ({10{received[351]}} & 10'b1011000110) ^ ({10{received[352]}} & 10'b0000110011) ^ ({10{received[353]}} & 10'b1100110000) ^ ({10{received[354]}} & 10'b1101101100) ^ ({10{received[355]}} & 10'b1010100101) ^ ({10{received[356]}} & 10'b1000001010) ^ ({10{received[357]}} & 10'b0011101000) ^ ({10{received[358]}} & 10'b1010011011) ^ ({10{received[359]}} & 10'b0111101010) ^ ({10{received[360]}} & 10'b1010011111) ^ ({10{received[361]}} & 10'b0110101010) ^ ({10{received[362]}} & 10'b1010010110) ^ ({10{received[363]}} & 10'b0100111010) ^ ({10{received[364]}} & 10'b1110000100) ^ ({10{received[365]}} & 10'b0000111110) ^ ({10{received[366]}} & 10'b1111100000) ^ ({10{received[367]}} & 10'b1001110111) ^ ({10{received[368]}} & 10'b1100110001) ^ ({10{received[369]}} & 10'b1101111100) ^ ({10{received[370]}} & 10'b1110100101) ^ ({10{received[371]}} & 10'b1000101110) ^ ({10{received[372]}} & 10'b1010101000) ^ ({10{received[373]}} & 10'b1011011010) ^ ({10{received[374]}} & 10'b0111110011) ^ ({10{received[375]}} & 10'b1100001111) ^ ({10{received[376]}} & 10'b0010011100) ^ ({10{received[377]}} & 10'b0111010010) ^ ({10{received[378]}} & 10'b0100011111) ^ ({10{received[379]}} & 10'b0111010100) ^ ({10{received[380]}} & 10'b0101111111) ^ ({10{received[381]}} & 10'b1111011101) ^ ({10{received[382]}} & 10'b0110100111) ^ ({10{received[383]}} & 10'b1001000110) ^ ({10{received[384]}} & 10'b0000100001) ^ ({10{received[385]}} & 10'b1000010000) ^ ({10{received[386]}} & 10'b0101001000) ^ ({10{received[387]}} & 10'b0010101101) ^ ({10{received[388]}} & 10'b1011000010) ^ ({10{received[389]}} & 10'b0001110011) ^ ({10{received[390]}} & 10'b1100111001) ^ ({10{received[391]}} & 10'b1111111100) ^ ({10{received[392]}} & 10'b1110110111) ^ ({10{received[393]}} & 10'b1100001110) ^ ({10{received[394]}} & 10'b0010001100) ^ ({10{received[395]}} & 10'b0011010010) ^ ({10{received[396]}} & 10'b0100111011) ^ ({10{received[397]}} & 10'b1110010100) ^ ({10{received[398]}} & 10'b0100111110) ^ ({10{received[399]}} & 10'b1111000100) ^ ({10{received[400]}} & 10'b0000110111) ^ ({10{received[401]}} & 10'b1101110000) ^ ({10{received[402]}} & 10'b1101100101) ^ ({10{received[403]}} & 10'b1000110101) ^ ({10{received[404]}} & 10'b1100011000) ^ ({10{received[405]}} & 10'b0111101100) ^ ({10{received[406]}} & 10'b1011111111) ^ ({10{received[407]}} & 10'b1110100011) ^ ({10{received[408]}} & 10'b1001001110) ^ ({10{received[409]}} & 10'b0010100001) ^ ({10{received[410]}} & 10'b1000000010) ^ ({10{received[411]}} & 10'b0001101000) ^ ({10{received[412]}} & 10'b1010001001) ^ ({10{received[413]}} & 10'b0011001010) ^ ({10{received[414]}} & 10'b0010111011) ^ ({10{received[415]}} & 10'b1110100010) ^ ({10{received[416]}} & 10'b1001011110) ^ ({10{received[417]}} & 10'b0110100001) ^ ({10{received[418]}} & 10'b1000100110) ^ ({10{received[419]}} & 10'b1000101000) ^ ({10{received[420]}} & 10'b1011001000) ^ ({10{received[421]}} & 10'b0011010011) ^ ({10{received[422]}} & 10'b0100101011) ^ ({10{received[423]}} & 10'b1010010100) ^ ({10{received[424]}} & 10'b0100011010) ^ ({10{received[425]}} & 10'b0110000100) ^ ({10{received[426]}} & 10'b0001110110) ^ ({10{received[427]}} & 10'b1101101001) ^ ({10{received[428]}} & 10'b1011110101) ^ ({10{received[429]}} & 10'b1100000011) ^ ({10{received[430]}} & 10'b0001011100) ^ ({10{received[431]}} & 10'b0111001001) ^ ({10{received[432]}} & 10'b0010101111) ^ ({10{received[433]}} & 10'b1011100010) ^ ({10{received[434]}} & 10'b1001110011) ^ ({10{received[435]}} & 10'b1101110001) ^ ({10{received[436]}} & 10'b1101110101) ^ ({10{received[437]}} & 10'b1100110101) ^ ({10{received[438]}} & 10'b1100111100) ^ ({10{received[439]}} & 10'b1110101100) ^ ({10{received[440]}} & 10'b1010111110) ^ ({10{received[441]}} & 10'b1110111010) ^ ({10{received[442]}} & 10'b1111011110) ^ ({10{received[443]}} & 10'b0110010111) ^ ({10{received[444]}} & 10'b0101000110) ^ ({10{received[445]}} & 10'b0001001101) ^ ({10{received[446]}} & 10'b0011011001) ^ ({10{received[447]}} & 10'b0110001011) ^ ({10{received[448]}} & 10'b0010000110) ^ ({10{received[449]}} & 10'b0001110010) ^ ({10{received[450]}} & 10'b1100101001) ^ ({10{received[451]}} & 10'b1011111100) ^ ({10{received[452]}} & 10'b1110010011) ^ ({10{received[453]}} & 10'b0101001110) ^ ({10{received[454]}} & 10'b0011001101) ^ ({10{received[455]}} & 10'b0011001011) ^ ({10{received[456]}} & 10'b0010101011) ^ ({10{received[457]}} & 10'b1010100010) ^ ({10{received[458]}} & 10'b1001111010) ^ ({10{received[459]}} & 10'b1111100001) ^ ({10{received[460]}} & 10'b1001100111) ^ ({10{received[461]}} & 10'b1000110001) ^ ({10{received[462]}} & 10'b1101011000) ^ ({10{received[463]}} & 10'b0111100101) ^ ({10{received[464]}} & 10'b1001101111) ^ ({10{received[465]}} & 10'b1010110001) ^ ({10{received[466]}} & 10'b1101001010) ^ ({10{received[467]}} & 10'b0011000101) ^ ({10{received[468]}} & 10'b0001001011) ^ ({10{received[469]}} & 10'b0010111001) ^ ({10{received[470]}} & 10'b1110000010) ^ ({10{received[471]}} & 10'b0001011110) ^ ({10{received[472]}} & 10'b0111101001) ^ ({10{received[473]}} & 10'b1010101111) ^ ({10{received[474]}} & 10'b1010101010) ^ ({10{received[475]}} & 10'b1011111010) ^ ({10{received[476]}} & 10'b1111110011) ^ ({10{received[477]}} & 10'b1101000111) ^ ({10{received[478]}} & 10'b0000010101) ^ ({10{received[479]}} & 10'b0101010000) ^ ({10{received[480]}} & 10'b0100101101) ^ ({10{received[481]}} & 10'b1011110100) ^ ({10{received[482]}} & 10'b1100010011) ^ ({10{received[483]}} & 10'b0101011100) ^ ({10{received[484]}} & 10'b0111101101) ^ ({10{received[485]}} & 10'b1011101111) ^ ({10{received[486]}} & 10'b1010100011) ^ ({10{received[487]}} & 10'b1001101010) ^ ({10{received[488]}} & 10'b1011100001) ^ ({10{received[489]}} & 10'b1001000011) ^ ({10{received[490]}} & 10'b0001110001) ^ ({10{received[491]}} & 10'b1100011001) ^ ({10{received[492]}} & 10'b0111111100) ^ ({10{received[493]}} & 10'b1111111111) ^ ({10{received[494]}} & 10'b1110000111) ^ ({10{received[495]}} & 10'b0000001110) ^ ({10{received[496]}} & 10'b0011100000) ^ ({10{received[497]}} & 10'b1000011011) ^ ({10{received[498]}} & 10'b0111111000) ^ ({10{received[499]}} & 10'b1110111111) ^ ({10{received[500]}} & 10'b1110001110) ^ ({10{received[501]}} & 10'b0010011110) ^ ({10{received[502]}} & 10'b0111110010) ^ ({10{received[503]}} & 10'b1100011111) ^ ({10{received[504]}} & 10'b0110011100) ^ ({10{received[505]}} & 10'b0111110110) ^ ({10{received[506]}} & 10'b1101011111) ^ ({10{received[507]}} & 10'b0110010101) ^ ({10{received[508]}} & 10'b0101100110) ^ ({10{received[509]}} & 10'b1001001101) ^ ({10{received[510]}} & 10'b0010010001) ^ ({10{received[511]}} & 10'b0100000010) ^ ({10{received[512]}} & 10'b0000000100) ^ ({10{received[513]}} & 10'b0001000000) ^ ({10{received[514]}} & 10'b0000001001) ^ ({10{received[515]}} & 10'b0010010000) ^ ({10{received[516]}} & 10'b0100010010) ^ ({10{received[517]}} & 10'b0100000100) ^ ({10{received[518]}} & 10'b0001100100) ^ ({10{received[519]}} & 10'b1001001001) ^ ({10{received[520]}} & 10'b0011010001) ^ ({10{received[521]}} & 10'b0100001011) ^ ({10{received[522]}} & 10'b0010010100) ^ ({10{received[523]}} & 10'b0101010010) ^ ({10{received[524]}} & 10'b0100001101) ^ ({10{received[525]}} & 10'b0011110100) ^ ({10{received[526]}} & 10'b1101011011) ^ ({10{received[527]}} & 10'b0111010101) ^ ({10{received[528]}} & 10'b0101101111) ^ ({10{received[529]}} & 10'b1011011101) ^ ({10{received[530]}} & 10'b0110000011) ^ ({10{received[531]}} & 10'b0000000110) ^ ({10{received[532]}} & 10'b0001100000) ^ ({10{received[533]}} & 10'b1000001001) ^ ({10{received[534]}} & 10'b0011011000) ^ ({10{received[535]}} & 10'b0110011011) ^ ({10{received[536]}} & 10'b0110000110) ^ ({10{received[537]}} & 10'b0001010110) ^ ({10{received[538]}} & 10'b0101101001) ^ ({10{received[539]}} & 10'b1010111101) ^ ({10{received[540]}} & 10'b1110001010) ^ ({10{received[541]}} & 10'b0011011110);
  assign syndrome5 = ({10{received[0]}} & 10'b0000000001) ^ 
  ({10{received[1]}} & 10'b0000100000) ^ ({10{received[2]}} & 10'b0000001001) ^ ({10{received[3]}} & 10'b0100100000) ^ ({10{received[4]}} & 10'b0001000001) ^ ({10{received[5]}} & 10'b0000110010) ^ ({10{received[6]}} & 10'b1001001001) ^ ({10{received[7]}} & 10'b0110100010) ^ ({10{received[8]}} & 10'b0000100101) ^ ({10{received[9]}} & 10'b0010101001) ^ ({10{received[10]}} & 10'b0100001101) ^ ({10{received[11]}} & 10'b0111101000) ^ ({10{received[12]}} & 10'b0101110111) ^ ({10{received[13]}} & 10'b1010110011) ^ ({10{received[14]}} & 10'b1011011101) ^ ({10{received[15]}} & 10'b1100000110) ^ ({10{received[16]}} & 10'b0000011000) ^ ({10{received[17]}} & 10'b1100000000) ^ ({10{received[18]}} & 10'b0011011000) ^ ({10{received[19]}} & 10'b1100110110) ^ ({10{received[20]}} & 10'b1000010001) ^ ({10{received[21]}} & 10'b1010110000) ^ ({10{received[22]}} & 10'b1010111101) ^ ({10{received[23]}} & 10'b1100011101) ^ ({10{received[24]}} & 10'b1101111000) ^ ({10{received[25]}} & 10'b1111000011) ^ ({10{received[26]}} & 10'b0010001110) ^ ({10{received[27]}} & 10'b0111100100) ^ ({10{received[28]}} & 10'b0011110111) ^ ({10{received[29]}} & 10'b1011011111) ^ ({10{received[30]}} & 10'b1101000110) ^ ({10{received[31]}} & 10'b0000001010) ^ ({10{received[32]}} & 10'b0101000000) ^ ({10{received[33]}} & 10'b0001011010) ^ ({10{received[34]}} & 10'b1101010010) ^ ({10{received[35]}} & 10'b1010001010) ^ ({10{received[36]}} & 10'b0111110100) ^ ({10{received[37]}} & 10'b1011110111) ^ ({10{received[38]}} & 10'b1001001111) ^ ({10{received[39]}} & 10'b0101100010) ^ ({10{received[40]}} & 10'b0000010011) ^ ({10{received[41]}} & 10'b1001100000) ^ ({10{received[42]}} & 10'b0010001011) ^ ({10{received[43]}} & 10'b0101000100) ^ ({10{received[44]}} & 10'b0011011010) ^ ({10{received[45]}} & 10'b1101110110) ^ ({10{received[46]}} & 10'b1000000011) ^ ({10{received[47]}} & 10'b0011110000) ^ ({10{received[48]}} & 10'b1000111111) ^ ({10{received[49]}} & 10'b1101111001) ^ ({10{received[50]}} & 10'b1111100011) ^ ({10{received[51]}} & 10'b0010000111) ^ ({10{received[52]}} & 10'b0011000100) ^ ({10{received[53]}} & 10'b0010110110) ^ ({10{received[54]}} & 10'b1011101101) ^ ({10{received[55]}} & 10'b0100001111) ^ ({10{received[56]}} & 10'b0110101000) ^ ({10{received[57]}} & 10'b0101100101) ^ ({10{received[58]}} & 10'b0011110011) ^ ({10{received[59]}} & 10'b1001011111) ^ ({10{received[60]}} & 10'b1101100010) ^ ({10{received[61]}} & 10'b0010000011) ^ ({10{received[62]}} & 10'b0001000100) ^ ({10{received[63]}} & 10'b0010010010) ^ ({10{received[64]}} & 10'b1001100100) ^ ({10{received[65]}} & 10'b0000001011) ^ ({10{received[66]}} & 10'b0101100000) ^ ({10{received[67]}} & 10'b0001010011) ^ ({10{received[68]}} & 10'b1001110010) ^ ({10{received[69]}} & 10'b1011001011) ^ ({10{received[70]}} & 10'b0111000110) ^ ({10{received[71]}} & 10'b0010111110) ^ ({10{received[72]}} & 10'b1111101101) ^ ({10{received[73]}} & 10'b0101000111) ^ ({10{received[74]}} & 10'b0010111010) ^ ({10{received[75]}} & 10'b1101101101) ^ ({10{received[76]}} & 10'b0101100011) ^ ({10{received[77]}} & 10'b0000110011) ^ ({10{received[78]}} & 10'b1001101001) ^ ({10{received[79]}} & 10'b0110101011) ^ ({10{received[80]}} & 10'b0100000101) ^ ({10{received[81]}} & 10'b0011101000) ^ ({10{received[82]}} & 10'b0100111111) ^ ({10{received[83]}} & 10'b1110100001) ^ ({10{received[84]}} & 10'b0011010101) ^ ({10{received[85]}} & 10'b1010010110) ^ ({10{received[86]}} & 10'b1001110100) ^ ({10{received[87]}} & 10'b1000001011) ^ ({10{received[88]}} & 10'b0111110000) ^ ({10{received[89]}} & 10'b1001110111) ^ ({10{received[90]}} & 10'b1001101011) ^ ({10{received[91]}} & 10'b0111101011) ^ ({10{received[92]}} & 10'b0100010111) ^ ({10{received[93]}} & 10'b1010101000) ^ ({10{received[94]}} & 10'b0110111101) ^ ({10{received[95]}} & 10'b1111000101) ^ ({10{received[96]}} & 10'b0001001110) ^ ({10{received[97]}} & 10'b0111010010) ^ ({10{received[98]}} & 10'b1000111110) ^ ({10{received[99]}} & 10'b1101011001) ^ ({10{received[100]}} & 10'b1111101010) ^ ({10{received[101]}} & 10'b0110100111) ^ ({10{received[102]}} & 10'b0010000101) ^ ({10{received[103]}} & 10'b0010000100) ^ ({10{received[104]}} & 10'b0010100100) ^ ({10{received[105]}} & 10'b0010101101) ^ ({10{received[106]}} & 10'b0110001101) ^ ({10{received[107]}} & 10'b0111001100) ^ ({10{received[108]}} & 10'b0111111110) ^ ({10{received[109]}} & 10'b1110110111) ^ ({10{received[110]}} & 10'b1000010101) ^ ({10{received[111]}} & 10'b1000110000) ^ ({10{received[112]}} & 10'b1010011001) ^ ({10{received[113]}} & 10'b1110010100) ^ ({10{received[114]}} & 10'b1001111100) ^ ({10{received[115]}} & 10'b1100001011) ^ ({10{received[116]}} & 10'b0110111000) ^ ({10{received[117]}} & 10'b1101100101) ^ ({10{received[118]}} & 10'b0001100011) ^ ({10{received[119]}} & 10'b0001111011) ^ ({10{received[120]}} & 10'b1101111011) ^ ({10{received[121]}} & 10'b1110100011) ^ ({10{received[122]}} & 10'b0010010101) ^ ({10{received[123]}} & 10'b1010000100) ^ ({10{received[124]}} & 10'b0000110100) ^ ({10{received[125]}} & 10'b1010001001) ^ ({10{received[126]}} & 10'b0110010100) ^ ({10{received[127]}} & 10'b1011101100) ^ ({10{received[128]}} & 10'b0100101111) ^ ({10{received[129]}} & 10'b0110100001) ^ ({10{received[130]}} & 10'b0001000101) ^ ({10{received[131]}} & 10'b0010110010) ^ ({10{received[132]}} & 10'b1001101101) ^ ({10{received[133]}} & 10'b0100101011) ^ ({10{received[134]}} & 10'b0100100001) ^ ({10{received[135]}} & 10'b0001100001) ^ ({10{received[136]}} & 10'b0000111011) ^ ({10{received[137]}} & 10'b1101101001) ^ ({10{received[138]}} & 10'b0111100011) ^ ({10{received[139]}} & 10'b0000010111) ^ ({10{received[140]}} & 10'b1011100000) ^ ({10{received[141]}} & 10'b0010101111) ^ ({10{received[142]}} & 10'b0111001101) ^ ({10{received[143]}} & 10'b0111011110) ^ ({10{received[144]}} & 10'b1110111110) ^ ({10{received[145]}} & 10'b1100110101) ^ ({10{received[146]}} & 10'b1001110001) ^ ({10{received[147]}} & 10'b1010101011) ^ ({10{received[148]}} & 10'b0111011101) ^ ({10{received[149]}} & 10'b1111011110) ^ ({10{received[150]}} & 10'b1100101110) ^ ({10{received[151]}} & 10'b0100010001) ^ ({10{received[152]}} & 10'b1001101000) ^ ({10{received[153]}} & 10'b0110001011) ^ ({10{received[154]}} & 10'b0100001100) ^ ({10{received[155]}} & 10'b0111001000) ^ ({10{received[156]}} & 10'b0101111110) ^ ({10{received[157]}} & 10'b1110010011) ^ ({10{received[158]}} & 10'b1010011100) ^ ({10{received[159]}} & 10'b1100110100) ^ ({10{received[160]}} & 10'b1001010001) ^ ({10{received[161]}} & 10'b1010100010) ^ ({10{received[162]}} & 10'b0011111101) ^ ({10{received[163]}} & 10'b1110011111) ^ ({10{received[164]}} & 10'b1100011100) ^ ({10{received[165]}} & 10'b1101011000) ^ ({10{received[166]}} & 10'b1111001010) ^ ({10{received[167]}} & 10'b0110101110) ^ ({10{received[168]}} & 10'b0110100101) ^ ({10{received[169]}} & 10'b0011000101) ^ ({10{received[170]}} & 10'b0010010110) ^ ({10{received[171]}} & 10'b1011100100) ^ ({10{received[172]}} & 10'b0000101111) ^ ({10{received[173]}} & 10'b0111101001) ^ ({10{received[174]}} & 10'b0101010111) ^ ({10{received[175]}} & 10'b1010111010) ^ ({10{received[176]}} & 10'b1111111101) ^ ({10{received[177]}} & 10'b1101000111) ^ ({10{received[178]}} & 10'b0000101010) ^ ({10{received[179]}} & 10'b0101001001) ^ ({10{received[180]}} & 10'b0101111010) ^ ({10{received[181]}} & 10'b1100010011) ^ ({10{received[182]}} & 10'b1010111000) ^ ({10{received[183]}} & 10'b1110111101) ^ ({10{received[184]}} & 10'b1101010101) ^ ({10{received[185]}} & 10'b1001101010) ^ ({10{received[186]}} & 10'b0111001011) ^ ({10{received[187]}} & 10'b0100011110) ^ ({10{received[188]}} & 10'b1110001000) ^ ({10{received[189]}} & 10'b0111111100) ^ ({10{received[190]}} & 10'b1111110111) ^ ({10{received[191]}} & 10'b1000000111) ^ ({10{received[192]}} & 10'b0001110000) ^ ({10{received[193]}} & 10'b1000011011) ^ ({10{received[194]}} & 10'b1111110000) ^ ({10{received[195]}} & 10'b1011100111) ^ ({10{received[196]}} & 10'b0001001111) ^ ({10{received[197]}} & 10'b0111110010) ^ ({10{received[198]}} & 10'b1000110111) ^ ({10{received[199]}} & 10'b1001111001) ^ ({10{received[200]}} & 10'b1110101011) ^ ({10{received[201]}} & 10'b0110010101) ^ ({10{received[202]}} & 10'b1011001100) ^ ({10{received[203]}} & 10'b0100100110) ^ ({10{received[204]}} & 10'b0010000001) ^ ({10{received[205]}} & 10'b0000000100) ^ ({10{received[206]}} & 10'b0010000000) ^ ({10{received[207]}} & 10'b0000100100) ^ ({10{received[208]}} & 10'b0010001001) ^ ({10{received[209]}} & 10'b0100000100) ^ ({10{received[210]}} & 10'b0011001000) ^ ({10{received[211]}} & 10'b0100110110) ^ ({10{received[212]}} & 10'b1010000001) ^ ({10{received[213]}} & 10'b0010010100) ^ ({10{received[214]}} & 10'b1010100100) ^ ({10{received[215]}} & 10'b0000111101) ^ ({10{received[216]}} & 10'b1110101001) ^ ({10{received[217]}} & 10'b0111010101) ^ ({10{received[218]}} & 10'b1011011110) ^ ({10{received[219]}} & 10'b1101100110) ^ ({10{received[220]}} & 10'b0000000011) ^ ({10{received[221]}} & 10'b0001100000) ^ ({10{received[222]}} & 10'b0000011011) ^ ({10{received[223]}} & 10'b1101100000) ^ ({10{received[224]}} & 10'b0011000011) ^ ({10{received[225]}} & 10'b0001010110) ^ ({10{received[226]}} & 10'b1011010010) ^ ({10{received[227]}} & 10'b1011100110) ^ ({10{received[228]}} & 10'b0001101111) ^ ({10{received[229]}} & 10'b0111111011) ^ ({10{received[230]}} & 10'b1100010111) ^ ({10{received[231]}} & 10'b1000111000) ^ ({10{received[232]}} & 10'b1110011001) ^ ({10{received[233]}} & 10'b1111011100) ^ ({10{received[234]}} & 10'b1101101110) ^ ({10{received[235]}} & 10'b0100000011) ^ ({10{received[236]}} & 10'b0000101000) ^ ({10{received[237]}} & 10'b0100001001) ^ ({10{received[238]}} & 10'b0101101000) ^ ({10{received[239]}} & 10'b0101010011) ^ ({10{received[240]}} & 10'b1000111010) ^ ({10{received[241]}} & 10'b1111011001) ^ ({10{received[242]}} & 10'b1111001110) ^ ({10{received[243]}} & 10'b0100101110) ^ ({10{received[244]}} & 10'b0110000001) ^ ({10{received[245]}} & 10'b0001001100) ^ ({10{received[246]}} & 10'b0110010010) ^ ({10{received[247]}} & 10'b1000101100) ^ ({10{received[248]}} & 10'b0100011001) ^ ({10{received[249]}} & 10'b1101101000) ^ ({10{received[250]}} & 10'b0111000011) ^ ({10{received[251]}} & 10'b0000011110) ^ ({10{received[252]}} & 10'b1111000000) ^ ({10{received[253]}} & 10'b0011101110) ^ ({10{received[254]}} & 10'b0111111111) ^ ({10{received[255]}} & 10'b1110010111) ^ ({10{received[256]}} & 10'b1000011100) ^ ({10{received[257]}} & 10'b1100010000) ^ ({10{received[258]}} & 10'b1011011000) ^ ({10{received[259]}} & 10'b1110100110) ^ ({10{received[260]}} & 10'b0000110101) ^ ({10{received[261]}} & 10'b1010101001) ^ ({10{received[262]}} & 10'b0110011101) ^ ({10{received[263]}} & 10'b1111001100) ^ ({10{received[264]}} & 10'b0101101110) ^ ({10{received[265]}} & 10'b0110010011) ^ ({10{received[266]}} & 10'b1000001100) ^ ({10{received[267]}} & 10'b0100010000) ^ ({10{received[268]}} & 10'b1001001000) ^ ({10{received[269]}} & 10'b0110000010) ^ ({10{received[270]}} & 10'b0000101100) ^ ({10{received[271]}} & 10'b0110001001) ^ ({10{received[272]}} & 10'b0101001100) ^ ({10{received[273]}} & 10'b0111011010) ^ ({10{received[274]}} & 10'b1100111110) ^ ({10{received[275]}} & 10'b1100010001) ^ ({10{received[276]}} & 10'b1011111000) ^ ({10{received[277]}} & 10'b1110101111) ^ ({10{received[278]}} & 10'b0100010101) ^ ({10{received[279]}} & 10'b1011101000) ^ ({10{received[280]}} & 10'b0110101111) ^ ({10{received[281]}} & 10'b0110000101) ^ ({10{received[282]}} & 10'b0011001100) ^ ({10{received[283]}} & 10'b0110110110) ^ ({10{received[284]}} & 10'b1010100101) ^ ({10{received[285]}} & 10'b0000011101) ^ ({10{received[286]}} & 10'b1110100000) ^ ({10{received[287]}} & 10'b0011110101) ^ ({10{received[288]}} & 10'b1010011111) ^ ({10{received[289]}} & 10'b1101010100) ^ ({10{received[290]}} & 10'b1001001010) ^ ({10{received[291]}} & 10'b0111000010) ^ ({10{received[292]}} & 10'b0000111110) ^ ({10{received[293]}} & 10'b1111001001) ^ ({10{received[294]}} & 10'b0111001110) ^ ({10{received[295]}} & 10'b0110111110) ^ ({10{received[296]}} & 10'b1110100101) ^ ({10{received[297]}} & 10'b0001010101) ^ ({10{received[298]}} & 10'b1010110010) ^ ({10{received[299]}} & 10'b1011111101) ^ ({10{received[300]}} & 10'b1100001111) ^ ({10{received[301]}} & 10'b0100111000) ^ ({10{received[302]}} & 10'b1101000001) ^ ({10{received[303]}} & 10'b0011101010) ^ ({10{received[304]}} & 10'b0101111111) ^ ({10{received[305]}} & 10'b1110110011) ^ ({10{received[306]}} & 10'b1010010101) ^ ({10{received[307]}} & 10'b1000010100) ^ ({10{received[308]}} & 10'b1000010000) ^ ({10{received[309]}} & 10'b1010010000) ^ ({10{received[310]}} & 10'b1010110100) ^ ({10{received[311]}} & 10'b1000111101) ^ ({10{received[312]}} & 10'b1100111001) ^ ({10{received[313]}} & 10'b1111110001) ^ ({10{received[314]}} & 10'b1011000111) ^ ({10{received[315]}} & 10'b0001000110) ^ ({10{received[316]}} & 10'b0011010010) ^ ({10{received[317]}} & 10'b1001110110) ^ ({10{received[318]}} & 10'b1001001011) ^ ({10{received[319]}} & 10'b0111100010) ^ ({10{received[320]}} & 10'b0000110111) ^ ({10{received[321]}} & 10'b1011101001) ^ ({10{received[322]}} & 10'b0110001111) ^ ({10{received[323]}} & 10'b0110001100) ^ ({10{received[324]}} & 10'b0111101100) ^ ({10{received[325]}} & 10'b0111110111) ^ ({10{received[326]}} & 10'b1010010111) ^ ({10{received[327]}} & 10'b1001010100) ^ ({10{received[328]}} & 10'b1000000010) ^ ({10{received[329]}} & 10'b0011010000) ^ ({10{received[330]}} & 10'b1000110110) ^ ({10{received[331]}} & 10'b1001011001) ^ ({10{received[332]}} & 10'b1110100010) ^ ({10{received[333]}} & 10'b0010110101) ^ ({10{received[334]}} & 10'b1010001101) ^ ({10{received[335]}} & 10'b0100010100) ^ ({10{received[336]}} & 10'b1011001000) ^ ({10{received[337]}} & 10'b0110100110) ^ ({10{received[338]}} & 10'b0010100101) ^ ({10{received[339]}} & 10'b0010001101) ^ ({10{received[340]}} & 10'b0110000100) ^ ({10{received[341]}} & 10'b0011101100) ^ ({10{received[342]}} & 10'b0110111111) ^ ({10{received[343]}} & 10'b1110000101) ^ ({10{received[344]}} & 10'b0001011100) ^ ({10{received[345]}} & 10'b1110010010) ^ ({10{received[346]}} & 10'b1010111100) ^ ({10{received[347]}} & 10'b1100111101) ^ ({10{received[348]}} & 10'b1101110001) ^ ({10{received[349]}} & 10'b1011100011) ^ ({10{received[350]}} & 10'b0011001111) ^ ({10{received[351]}} & 10'b0111010110) ^ ({10{received[352]}} & 10'b1010111110) ^ ({10{received[353]}} & 10'b1101111101) ^ ({10{received[354]}} & 10'b1101100011) ^ ({10{received[355]}} & 10'b0010100011) ^ ({10{received[356]}} & 10'b0001001101) ^ ({10{received[357]}} & 10'b0110110010) ^ ({10{received[358]}} & 10'b1000100101) ^ ({10{received[359]}} & 10'b0000111001) ^ ({10{received[360]}} & 10'b1100101001) ^ ({10{received[361]}} & 10'b0111110001) ^ ({10{received[362]}} & 10'b1001010111) ^ ({10{received[363]}} & 10'b1001100010) ^ ({10{received[364]}} & 10'b0011001011) ^ ({10{received[365]}} & 10'b0101010110) ^ ({10{received[366]}} & 10'b1010011010) ^ ({10{received[367]}} & 10'b1111110100) ^ ({10{received[368]}} & 10'b1001100111) ^ ({10{received[369]}} & 10'b0001101011) ^ ({10{received[370]}} & 10'b0101111011) ^ ({10{received[371]}} & 10'b1100110011) ^ ({10{received[372]}} & 10'b1010110001) ^ ({10{received[373]}} & 10'b1010011101) ^ ({10{received[374]}} & 10'b1100010100) ^ ({10{received[375]}} & 10'b1001011000) ^ ({10{received[376]}} & 10'b1110000010) ^ ({10{received[377]}} & 10'b0010111100) ^ ({10{received[378]}} & 10'b1110101101) ^ ({10{received[379]}} & 10'b0101010101) ^ ({10{received[380]}} & 10'b1011111010) ^ ({10{received[381]}} & 10'b1111101111) ^ ({10{received[382]}} & 10'b0100000111) ^ ({10{received[383]}} & 10'b0010101000) ^ ({10{received[384]}} & 10'b0100101101) ^ ({10{received[385]}} & 10'b0111100001) ^ ({10{received[386]}} & 10'b0001010111) ^ ({10{received[387]}} & 10'b1011110010) ^ ({10{received[388]}} & 10'b1011101111) ^ ({10{received[389]}} & 10'b0101001111) ^ ({10{received[390]}} & 10'b0110111010) ^ ({10{received[391]}} & 10'b1100100101) ^ ({10{received[392]}} & 10'b0001110001) ^ ({10{received[393]}} & 10'b1000111011) ^ ({10{received[394]}} & 10'b1111111001) ^ ({10{received[395]}} & 10'b1111000111) ^ ({10{received[396]}} & 10'b0000001110) ^ ({10{received[397]}} & 10'b0111000000) ^ ({10{received[398]}} & 10'b0001111110) ^ ({10{received[399]}} & 10'b1111011011) ^ ({10{received[400]}} & 10'b1110001110) ^ ({10{received[401]}} & 10'b0100111100) ^ ({10{received[402]}} & 10'b1111000001) ^ ({10{received[403]}} & 10'b0011001110) ^ ({10{received[404]}} & 10'b0111110110) ^ ({10{received[405]}} & 10'b1010110111) ^ ({10{received[406]}} & 10'b1001011101) ^ ({10{received[407]}} & 10'b1100100010) ^ ({10{received[408]}} & 10'b0010010001) ^ ({10{received[409]}} & 10'b1000000100) ^ ({10{received[410]}} & 10'b0000010000) ^ ({10{received[411]}} & 10'b1000000000) ^ ({10{received[412]}} & 10'b0010010000) ^ ({10{received[413]}} & 10'b1000100100) ^ ({10{received[414]}} & 10'b0000011001) ^ ({10{received[415]}} & 10'b1100100000) ^ ({10{received[416]}} & 10'b0011010001) ^ ({10{received[417]}} & 10'b1000010110) ^ ({10{received[418]}} & 10'b1001010000) ^ ({10{received[419]}} & 10'b1010000010) ^ ({10{received[420]}} & 10'b0011110100) ^ ({10{received[421]}} & 10'b1010111111) ^ ({10{received[422]}} & 10'b1101011101) ^ ({10{received[423]}} & 10'b1101101010) ^ ({10{received[424]}} & 10'b0110000011) ^ ({10{received[425]}} & 10'b0000001100) ^ ({10{received[426]}} & 10'b0110000000) ^ ({10{received[427]}} & 10'b0001101100) ^ ({10{received[428]}} & 10'b0110011011) ^ ({10{received[429]}} & 10'b1100001100) ^ ({10{received[430]}} & 10'b0101011000) ^ ({10{received[431]}} & 10'b1101011010) ^ ({10{received[432]}} & 10'b1110001010) ^ ({10{received[433]}} & 10'b0110111100) ^ ({10{received[434]}} & 10'b1111100101) ^ ({10{received[435]}} & 10'b0001000111) ^ ({10{received[436]}} & 10'b0011110010) ^ ({10{received[437]}} & 10'b1001111111) ^ ({10{received[438]}} & 10'b1101101011) ^ ({10{received[439]}} & 10'b0110100011) ^ ({10{received[440]}} & 10'b0000000101) ^ ({10{received[441]}} & 10'b0010100000) ^ ({10{received[442]}} & 10'b0000101101) ^ ({10{received[443]}} & 10'b0110101001) ^ ({10{received[444]}} & 10'b0101000101) ^ ({10{received[445]}} & 10'b0011111010) ^ ({10{received[446]}} & 10'b1101111111) ^ ({10{received[447]}} & 10'b1100100011) ^ ({10{received[448]}} & 10'b0010110001) ^ ({10{received[449]}} & 10'b1000001101) ^ ({10{received[450]}} & 10'b0100110000) ^ ({10{received[451]}} & 10'b1001000001) ^ ({10{received[452]}} & 10'b0010100010) ^ ({10{received[453]}} & 10'b0001101101) ^ ({10{received[454]}} & 10'b0110111011) ^ ({10{received[455]}} & 10'b1100000101) ^ ({10{received[456]}} & 10'b0001111000) ^ ({10{received[457]}} & 10'b1100011011) ^ ({10{received[458]}} & 10'b1110111000) ^ ({10{received[459]}} & 10'b1111110101) ^ ({10{received[460]}} & 10'b1001000111) ^ ({10{received[461]}} & 10'b0001100010) ^ ({10{received[462]}} & 10'b0001011011) ^ ({10{received[463]}} & 10'b1101110010) ^ ({10{received[464]}} & 10'b1010000011) ^ ({10{received[465]}} & 10'b0011010100) ^ ({10{received[466]}} & 10'b1010110110) ^ ({10{received[467]}} & 10'b1001111101) ^ ({10{received[468]}} & 10'b1100101011) ^ ({10{received[469]}} & 10'b0110110001) ^ ({10{received[470]}} & 10'b1001000101) ^ ({10{received[471]}} & 10'b0000100010) ^ ({10{received[472]}} & 10'b0001001001) ^ ({10{received[473]}} & 10'b0100110010) ^ ({10{received[474]}} & 10'b1000000001) ^ ({10{received[475]}} & 10'b0010110000) ^ ({10{received[476]}} & 10'b1000101101) ^ ({10{received[477]}} & 10'b0100111001) ^ ({10{received[478]}} & 10'b1101100001) ^ ({10{received[479]}} & 10'b0011100011) ^ ({10{received[480]}} & 10'b0001011111) ^ ({10{received[481]}} & 10'b1111110010) ^ ({10{received[482]}} & 10'b1010100111) ^ ({10{received[483]}} & 10'b0001011101) ^ ({10{received[484]}} & 10'b1110110010) ^ ({10{received[485]}} & 10'b1010110101) ^ ({10{received[486]}} & 10'b1000011101) ^ ({10{received[487]}} & 10'b1100110000) ^ ({10{received[488]}} & 10'b1011010001) ^ ({10{received[489]}} & 10'b1010000110) ^ ({10{received[490]}} & 10'b0001110100) ^ ({10{received[491]}} & 10'b1010011011) ^ ({10{received[492]}} & 10'b1111010100) ^ ({10{received[493]}} & 10'b1001101110) ^ ({10{received[494]}} & 10'b0101001011) ^ ({10{received[495]}} & 10'b0100111010) ^ ({10{received[496]}} & 10'b1100000001) ^ ({10{received[497]}} & 10'b0011111000) ^ ({10{received[498]}} & 10'b1100111111) ^ ({10{received[499]}} & 10'b1100110001) ^ ({10{received[500]}} & 10'b1011110001) ^ ({10{received[501]}} & 10'b1010001111) ^ ({10{received[502]}} & 10'b0101010100) ^ ({10{received[503]}} & 10'b1011011010) ^ ({10{received[504]}} & 10'b1111100110) ^ ({10{received[505]}} & 10'b0000100111) ^ ({10{received[506]}} & 10'b0011101001) ^ ({10{received[507]}} & 10'b0100011111) ^ ({10{received[508]}} & 10'b1110101000) ^ ({10{received[509]}} & 10'b0111110101) ^ ({10{received[510]}} & 10'b1011010111) ^ ({10{received[511]}} & 10'b1001000110) ^ ({10{received[512]}} & 10'b0001000010) ^ ({10{received[513]}} & 10'b0001010010) ^ ({10{received[514]}} & 10'b1001010010) ^ ({10{received[515]}} & 10'b1011000010) ^ ({10{received[516]}} & 10'b0011100110) ^ ({10{received[517]}} & 10'b0011111111) ^ ({10{received[518]}} & 10'b1111011111) ^ ({10{received[519]}} & 10'b1100001110) ^ ({10{received[520]}} & 10'b0100011000) ^ ({10{received[521]}} & 10'b1101001000) ^ ({10{received[522]}} & 10'b0111001010) ^ ({10{received[523]}} & 10'b0100111110) ^ ({10{received[524]}} & 10'b1110000001) ^ ({10{received[525]}} & 10'b0011011100) ^ ({10{received[526]}} & 10'b1110110110) ^ ({10{received[527]}} & 10'b1000110101) ^ ({10{received[528]}} & 10'b1000111001) ^ ({10{received[529]}} & 10'b1110111001) ^ ({10{received[530]}} & 10'b1111010101) ^ ({10{received[531]}} & 10'b1001001110) ^ ({10{received[532]}} & 10'b0101000010) ^ ({10{received[533]}} & 10'b0000011010) ^ ({10{received[534]}} & 10'b1101000000) ^ ({10{received[535]}} & 10'b0011001010) ^ ({10{received[536]}} & 10'b0101110110) ^ ({10{received[537]}} & 10'b1010010011) ^ ({10{received[538]}} & 10'b1011010100) ^ ({10{received[539]}} & 10'b1000100110) ^ ({10{received[540]}} & 10'b0001011001) ^ ({10{received[541]}} & 10'b1100110010);
endmodule