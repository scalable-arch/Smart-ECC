module SEC_encoder(input [127:0] message, output [135:0] codeword);

	assign codeword[135:8] = message[127:0];
	assign codeword[7] = ^(message&128'b10101010011110000110010100100110001101110110110001010101011110100111001011010111110111111111100010110101011001010000101101100110);
	assign codeword[6] = ^(message&128'b01001101100111000100011011100010101110001100101110110111011001101110001100001100011110011100001001111001001101111001010010001110);
	assign codeword[5] = ^(message&128'b10010000100100101010111111101101001111111111001101100101110000111001010010111001011110001011010010101001100100011010011100100011);
	assign codeword[4] = ^(message&128'b00010111111101011111111001100000000000100000110011000011010000011011010100011011101000010100110110111010001010110111110101110111);
	assign codeword[3] = ^(message&128'b11010101011000000010101010011011110100101111001110000011111010110110110010010000101001101010000100011111011001010100110111011110);
	assign codeword[2] = ^(message&128'b00011000010000010100010011010101100000111110000010111110111111010001100111111010100111011000111110101100101011011011111000111100);
	assign codeword[1] = ^(message&128'b11101100001010110011110110100100010010110011111000101110101111111110100100001111111100111000010011001001101000110100000000011011);
	assign codeword[0] = ^(message&128'b10111110011111101101111001011000010100111000101010101000110010101101001111100011010111001001011001011010011111000000000110011010);

endmodule
